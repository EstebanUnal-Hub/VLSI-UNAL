* Generated from tt_um_mult_4.tim
* VDD Level: 3.3 V

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.tran 1e-11 1.32e-06
.print tran format=raw file=tt_um_mult_4.raw v(*)

* Power rails
Vvdd VPWR 0 DC 3.3
Vgnd VGND 0 DC 0

* clk
V_clk clk 0 PWL(0 0 9.999e-09 0 1e-08 3.3 1.9999e-08 3.3 2e-08 0 2.9999e-08 0 3e-08 3.3 3.9999e-08 3.3 4e-08 0 4.9999e-08 0 5e-08 3.3 5.9999e-08 3.3 6e-08 0 6.9999e-08 0 7e-08 3.3 7.9999e-08 3.3 8e-08 0 8.9999e-08 0 9e-08 3.3 9.9999e-08 3.3 1e-07 0 1.09999e-07 0 1.1e-07 3.3 1.19999e-07 3.3 1.2e-07 0 1.29999e-07 0 1.3e-07 3.3 1.39999e-07 3.3 1.4e-07 0 1.49999e-07 0 1.5e-07 3.3 1.59999e-07 3.3 1.6e-07 0 1.69999e-07 0 1.7e-07 3.3 1.79999e-07 3.3 1.8e-07 0 1.89999e-07 0 1.9e-07 3.3 1.99999e-07 3.3 2e-07 0 2.09999e-07 0 2.1e-07 3.3 2.19999e-07 3.3 2.2e-07 0 2.29999e-07 0 2.3e-07 3.3 2.39999e-07 3.3 2.4e-07 0 2.49999e-07 0 2.5e-07 3.3 2.59999e-07 3.3 2.6e-07 0 2.69999e-07 0 2.7e-07 3.3 2.79999e-07 3.3 2.8e-07 0 2.89999e-07 0 2.9e-07 3.3 2.99999e-07 3.3 3e-07 0 3.09999e-07 0 3.1e-07 3.3 3.19999e-07 3.3 3.2e-07 0 3.29999e-07 0 3.3e-07 3.3 3.39999e-07 3.3 3.4e-07 0 3.49999e-07 0 3.5e-07 3.3 3.59999e-07 3.3 3.6e-07 0 3.69999e-07 0 3.7e-07 3.3 3.79999e-07 3.3 3.8e-07 0 3.89999e-07 0 3.9e-07 3.3 3.99999e-07 3.3 4e-07 0 4.09999e-07 0 4.1e-07 3.3 4.19999e-07 3.3 4.2e-07 0 4.29999e-07 0 4.3e-07 3.3 4.39999e-07 3.3 4.4e-07 0 4.49999e-07 0 4.5e-07 3.3 4.59999e-07 3.3 4.6e-07 0 4.69999e-07 0 4.7e-07 3.3 4.79999e-07 3.3 4.8e-07 0 4.89999e-07 0 4.9e-07 3.3 4.99999e-07 3.3 5e-07 0 5.09999e-07 0 5.1e-07 3.3 5.19999e-07 3.3 5.2e-07 0 5.29999e-07 0 5.3e-07 3.3 5.39999e-07 3.3 5.4e-07 0 5.49999e-07 0 5.5e-07 3.3 5.59999e-07 3.3 5.6e-07 0 5.69999e-07 0 5.7e-07 3.3 5.79999e-07 3.3 5.8e-07 0 5.89999e-07 0 5.9e-07 3.3 5.99999e-07 3.3 6e-07 0 6.09999e-07 0 6.1e-07 3.3 6.19999e-07 3.3 6.2e-07 0 6.29999e-07 0 6.3e-07 3.3 6.39999e-07 3.3 6.4e-07 0 6.49999e-07 0 6.5e-07 3.3 6.59999e-07 3.3 6.6e-07 0 6.69999e-07 0 6.7e-07 3.3 6.79999e-07 3.3 6.8e-07 0 6.89999e-07 0 6.9e-07 3.3 6.99999e-07 3.3 7e-07 0 7.09999e-07 0 7.1e-07 3.3 7.19999e-07 3.3 7.2e-07 0 7.29999e-07 0 7.3e-07 3.3 7.39999e-07 3.3 7.4e-07 0 7.49999e-07 0 7.5e-07 3.3 7.59999e-07 3.3 7.6e-07 0 7.69999e-07 0 7.7e-07 3.3 7.79999e-07 3.3 7.8e-07 0 7.89999e-07 0 7.9e-07 3.3 7.99999e-07 3.3 8e-07 0 8.09999e-07 0 8.1e-07 3.3 8.19999e-07 3.3 8.2e-07 0 8.29999e-07 0 8.3e-07 3.3 8.39999e-07 3.3 8.4e-07 0 8.49999e-07 0 8.5e-07 3.3 8.59999e-07 3.3 8.6e-07 0 8.69999e-07 0 8.7e-07 3.3 8.79999e-07 3.3 8.8e-07 0 8.89999e-07 0 8.9e-07 3.3 8.99999e-07 3.3 9e-07 0 9.09999e-07 0 9.1e-07 3.3 9.19999e-07 3.3 9.2e-07 0 9.29999e-07 0 9.3e-07 3.3 9.39999e-07 3.3 9.4e-07 0 9.49999e-07 0 9.5e-07 3.3 9.59999e-07 3.3 9.6e-07 0 9.69999e-07 0 9.7e-07 3.3 9.79999e-07 3.3 9.8e-07 0 9.89999e-07 0 9.9e-07 3.3 9.99999e-07 3.3 1e-06 0 1.009999e-06 0 1.01e-06 3.3 1.019999e-06 3.3 1.02e-06 0 1.029999e-06 0 1.03e-06 3.3 1.039999e-06 3.3 1.04e-06 0 1.049999e-06 0 1.05e-06 3.3 1.059999e-06 3.3 1.06e-06 0 1.069999e-06 0 1.07e-06 3.3 1.079999e-06 3.3 1.08e-06 0 1.089999e-06 0 1.09e-06 3.3 1.099999e-06 3.3 1.1e-06 0 1.109999e-06 0 1.11e-06 3.3 1.119999e-06 3.3 1.12e-06 0 1.129999e-06 0 1.13e-06 3.3 1.139999e-06 3.3 1.14e-06 0 1.149999e-06 0 1.15e-06 3.3 1.159999e-06 3.3 1.16e-06 0 1.169999e-06 0 1.17e-06 3.3 1.179999e-06 3.3 1.18e-06 0 1.189999e-06 0 1.19e-06 3.3 1.199999e-06 3.3 1.2e-06 0)

* done
V_done done 0 PWL(0 0 3.69999e-07 0 3.7e-07 3.3 5.69999e-07 3.3 5.7e-07 0)

* rst_n
V_rst_n rst_n 0 PWL(0 3.3 3.9999e-08 3.3 4e-08 0)

* ui_in[0]
V_ui_in[0] ui_in[0] 0 PWL(0 3.3)

* ui_in[1]
V_ui_in[1] ui_in[1] 0 PWL(0 0)

* ui_in[2]
V_ui_in[2] ui_in[2] 0 PWL(0 3.3)

* ui_in[3]
V_ui_in[3] ui_in[3] 0 PWL(0 0)

* ui_in[4]
V_ui_in[4] ui_in[4] 0 PWL(0 3.3)

* ui_in[5]
V_ui_in[5] ui_in[5] 0 PWL(0 0)

* ui_in[6]
V_ui_in[6] ui_in[6] 0 PWL(0 3.3)

* ui_in[7]
V_ui_in[7] ui_in[7] 0 PWL(0 3.3)

* uio_in[0]
V_uio_in[0] uio_in[0] 0 PWL(0 0 6.9999e-08 0 7e-08 3.3 1.09999e-07 3.3 1.1e-07 0)

.include "./tt_um_mult_4.spice"
.end
