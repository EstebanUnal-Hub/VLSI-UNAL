* NGSPICE file created from tt_um_femto.ext - technology: sky130A

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VNB VPB VGND VPWR X A1 A2 B1 C1
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10563 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10187 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB X A
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 VNB VPB VPWR VGND X S A1 A0
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.10887 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.27463 pd=1.495 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.27463 ps=1.495 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10887 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VNB VPB VGND VPWR X A2 A1 B1_N
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25837 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25837 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VPB VNB VGND VPWR
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X20 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09912 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 VNB VPB VPWR VGND A_N X B
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10187 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.07438 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10238 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10238 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VPB VNB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_4 VNB VPB VGND VPWR X C1 B1 A2 A1
X0 VGND A1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.104 ps=0.97 w=0.65 l=0.15
X1 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A1 a_1122_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2525 pd=1.505 as=0.14 ps=1.28 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2525 ps=1.505 w=1 l=0.15
X8 a_950_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X9 a_557_47# B1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 a_474_47# B1 a_748_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X11 VGND A2 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_79_21# C1 a_557_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14462 pd=1.095 as=0.06825 ps=0.86 w=0.65 l=0.15
X15 a_474_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X17 a_748_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.14462 ps=1.095 w=0.65 l=0.15
X18 a_474_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X19 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.195 ps=1.39 w=1 l=0.15
X20 a_79_21# A2 a_950_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 a_1122_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 VNB VPB VGND VPWR X D_N C B A
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 VNB VPB VGND VPWR X A2 A1 B1 C1
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11537 pd=1.005 as=0.13325 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.19987 pd=1.265 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.19987 ps=1.265 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.11537 ps=1.005 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd1_1 VPWR VGND VPB VNB X A
X0 X a_299_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1 VPWR a_193_47# a_299_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 VGND a_193_47# a_299_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X a_299_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VPB VNB VGND VPWR C B A Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_2 VPB VNB VGND VPWR A B C Y
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A1 A2 A3 B1 VPB VNB VGND VPWR
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VNB VPB VPWR VGND X A1_N A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.09862 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.09862 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VPB VNB VGND VPWR A_N B Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.09912 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_4 VNB VPB VGND VPWR B1 B2 A2_N A1_N X
X0 a_27_47# a_415_21# a_193_297# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_415_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3 a_415_21# A2_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_193_297# a_415_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_717_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_717_47# A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_27_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A1_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_193_297# a_415_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR a_415_21# a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X23 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_415_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VGND B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VNB VPB VGND VPWR B1_N A1 A2 X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPB VNB VPWR VGND X A1 A2 A3 B2 B1
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VPB VNB VGND VPWR Y B C A_N
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12513 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12513 ps=1.035 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_4 VNB VPB VGND VPWR C_N X A B
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.16737 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.16737 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.1312 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1778 pd=1.415 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1312 pd=1.05 as=0.2288 ps=1.355 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.05775 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2288 pd=1.355 as=0.1778 ps=1.415 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17325 pd=1.245 as=0.06825 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.17325 ps=1.245 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1728 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 VNB VPB VGND VPWR A_N B_N C D X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPB VNB VPWR VGND A1 B1_N Y A2
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VPB VNB VGND VPWR A1 A2 B1 B2 Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11537 ps=1.005 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.11537 pd=1.005 as=0.09262 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2325 ps=1.465 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2325 pd=1.465 as=0.1125 ps=1.225 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1125 pd=1.225 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09262 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_1 VPB VNB Y C1 B1 A1 A2 A3 VPWR VGND
X0 Y A1 a_194_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11537 pd=1.005 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_194_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X2 Y C1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1725 ps=1.345 w=1 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11213 ps=0.995 w=0.65 l=0.15
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.11537 ps=1.005 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7 a_376_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.165 ps=1.33 w=1 l=0.15
X8 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_12 VPB VNB VGND VPWR A X
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.135 ps=1.27 w=1 l=0.15
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10187 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 VNB VPB VGND VPWR A2 B1 Y A1
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR VNB VPB Q D CLK
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09262 ps=0.935 w=0.65 l=0.15
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10563 ps=0.975 w=0.65 l=0.15
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.09262 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X25 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X26 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_4 VNB VPB VGND VPWR B1_N X A2 A1
X0 VPWR B1_N a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.38 ps=2.76 w=1 l=0.15
X1 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3 a_575_47# a_27_297# a_187_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_743_297# A2 a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_27_297# a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_187_21# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_187_21# a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_187_21# a_27_297# a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VGND B1_N a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.91 w=0.65 l=0.15
X10 VGND A2 a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A1 a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_575_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_575_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 VNB VPB VGND VPWR A_N Y B
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 VPB VNB VPWR VGND B C A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_16 Y A VGND VPWR VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.2175 ps=1.435 w=1 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.275 ps=2.55 w=1 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.1575 ps=1.315 w=1 l=0.15
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09135 pd=0.855 as=0.06615 ps=0.735 w=0.42 l=0.15
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.09135 ps=0.855 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_4 VNB VPB VGND VPWR X B2 A1 A2 B1
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VPB VNB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_2 VPWR VGND VPB VNB B2 B1 A1 A2 X
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10238 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10238 ps=0.965 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1575 ps=1.315 w=1 l=0.15
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_4 VNB VPB VGND VPWR A3 A2 A1 B1 Y B2
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3375 pd=1.675 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2525 pd=1.505 as=0.3375 ps=1.675 w=1 l=0.15
X12 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X16 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13325 ps=1.06 w=0.65 l=0.15
X23 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2525 ps=1.505 w=1 l=0.15
X28 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X30 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 VPWR VGND VPB VNB C D_N X A B
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16835 pd=1.495 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1693 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.16835 ps=1.495 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1693 pd=1.5 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.10025 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB Y C1 B1 A1 A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VPB VNB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19627 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.19627 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_4 VGND VPWR VPB VNB X A2 A1 A3 B1
X0 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X8 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X10 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X14 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X15 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X18 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.145 ps=1.29 w=1 l=0.15
X22 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 VPB VNB VGND VPWR A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10187 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_2 VNB VPB VPWR VGND A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinvlp_4 VNB VPB VPWR VGND A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 VGND A a_268_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X3 Y A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X5 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X6 a_268_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
.ends

.subckt sky130_fd_sc_hd__inv_6 VPB VNB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_4 VNB VPB VGND VPWR A1 A2 B2 Y B1
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 VPB VNB VGND VPWR Y B A
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VNB VPB VGND VPWR A2 A1 Y B1
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_4 VNB VPB VGND VPWR A2 A1 C1 X B1
X0 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X3 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X4 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0.10887 pd=0.985 as=0.104 ps=0.97 w=0.65 l=0.15
X5 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.09262 ps=0.935 w=0.65 l=0.15
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X7 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X8 a_473_297# B1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16 ps=1.32 w=1 l=0.15
X9 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.12675 ps=1.04 w=0.65 l=0.15
X11 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10887 ps=0.985 w=0.65 l=0.15
X12 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0.09262 pd=0.935 as=0.09588 ps=0.945 w=0.65 l=0.15
X13 a_1123_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_555_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X15 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X16 VGND A2 a_1123_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.091 ps=0.93 w=0.65 l=0.15
X17 a_951_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.13975 ps=1.08 w=0.65 l=0.15
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X20 a_79_204# A1 a_951_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 a_79_204# C1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 a_727_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X23 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10187 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_4 VNB VPB VGND VPWR B A X
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11537 ps=1.005 w=0.65 l=0.15
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11537 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_2 VNB VPB VGND VPWR A_N X C D B_N
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.33075 ps=1.705 w=0.42 l=0.15
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33075 pd=1.705 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 X A1 A2 A3 B1 C1 VPB VNB VGND VPWR
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.11863 ps=1.015 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.20312 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.20312 ps=1.275 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_12 VNB VPB VGND VPWR Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.515 pd=3.03 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.33475 pd=2.33 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_16 VPB VNB VGND VPWR Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 VGND VPWR C A_N X D B VPB VNB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_4 VNB VPB VPWR VGND D C B A X
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__bufinv_8 VNB VPB VGND VPWR A Y
X0 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND a_215_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR a_215_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X22 Y a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_2 VPWR VGND VPB VNB X A1 A2 A3 B1 C1
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.20312 ps=1.275 w=0.65 l=0.15
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.20312 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.11863 ps=1.015 w=0.65 l=0.15
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_4 VNB VPB VGND VPWR B A X C_N D_N
X0 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2 a_315_380# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR A a_583_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_410# a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X7 a_583_297# B a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_315_380# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_397_297# a_205_93# a_315_380# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.25793 ps=2.52 w=1 l=0.15
X10 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X11 X a_315_380# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_499_297# a_27_410# a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X13 VPWR a_315_380# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X15 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11295 pd=1.4 as=0.1226 ps=1.32 w=0.42 l=0.15
X16 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND a_315_380# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_315_380# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X19 X a_315_380# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_2 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_1 VPB VNB VPWR VGND A C D Y B
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 VNB VPB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13487 ps=1.065 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12513 pd=1.035 as=0.11213 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.12513 ps=1.035 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.13487 pd=1.065 as=0.10563 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_4 VNB VPB VGND VPWR A_N C D X B_N
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_174_21# a_832_21# a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_832_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1764 ps=1.68 w=0.42 l=0.15
X4 a_766_47# a_27_47# a_652_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1365 ps=1.07 w=0.65 l=0.15
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_652_47# C a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 a_832_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.31165 ps=2.125 w=0.42 l=0.15
X10 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X11 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_556_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.11375 ps=1 w=0.65 l=0.15
X13 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.175 ps=1.35 w=1 l=0.15
X14 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR a_832_21# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31165 pd=2.125 as=0.165 ps=1.33 w=1 l=0.15
X18 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.21 ps=1.42 w=1 l=0.15
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_8 VNB VPB VGND VPWR A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1375 ps=1.275 w=1 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10187 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 VNB VPB VGND VPWR Y B A
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 VNB VPB VGND VPWR X D C B A
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_2 VPB VNB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.13975 pd=1.08 as=0.13325 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.1105 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12025 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13975 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_4 VNB VPB VGND VPWR B2 Y A2 A1 B1 C1
X0 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X10 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X14 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X26 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X32 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_8 VNB VPB VGND VPWR Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_4 VNB VPB VPWR VGND A2 A1 X B1
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 VNB VPB VPWR VGND A Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1659 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1386 ps=1.5 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_4 VPB VNB VGND VPWR B Y A
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VNB VPB VPWR VGND X D1 C1 B1 A2 A1
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.2125 ps=1.425 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.11863 ps=1.015 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.19825 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.19825 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.2175 ps=1.435 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.11863 ps=1.015 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3825 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2175 pd=1.435 as=0.3825 ps=1.765 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10563 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_4 VNB VPB VGND VPWR A X B
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.13813 ps=1.075 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13813 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB B1_N Y A1 A2
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10187 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_4 VNB VPB VGND VPWR A1 B1 B2 A2 X
X0 VPWR B1 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_484_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_566_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_96_21# B2 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A1 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 a_484_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_566_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X13 a_484_47# B2 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_96_21# A2 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_918_297# A2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_484_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_918_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_96_21# B1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 VGND A2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_96_21# B2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 VNB VPB VPWR VGND B1 Y A1 A2
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41ai_2 VNB VPB VGND VPWR A1 A2 A3 A4 Y B1
X0 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X4 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_299_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_549_297# A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_299_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A4 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_743_297# A2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_549_297# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 VPB VNB VGND VPWR X B1 A4 A3 A2 A1
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_1 VPB VNB VGND VPWR D_N C Y B A
X0 Y a_91_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_91_199# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_341_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X6 a_245_297# C a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_341_297# B a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X8 a_91_199# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X9 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.52 ps=3.04 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtn_1 VGND VPWR VPB VNB Q D GATE_N
X0 VPWR D a_299_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1 a_560_47# a_27_47# a_465_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.054 pd=0.66 as=0.066 ps=0.745 w=0.36 l=0.15
X2 a_465_47# a_299_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR GATE_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 VGND a_560_47# a_715_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR a_560_47# a_715_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X7 a_650_47# a_193_47# a_560_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.054 ps=0.66 w=0.36 l=0.15
X8 Q a_715_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X9 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X10 VPWR a_715_21# a_644_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 VGND D a_299_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 Q a_715_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X13 a_644_413# a_27_47# a_560_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_465_369# a_299_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_560_47# a_193_47# a_465_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X16 VGND GATE_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND a_715_21# a_650_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 VGND VPWR VPB VNB X A1 A2 A3 B1
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.26325 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.2125 ps=1.425 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.11375 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_4 VNB VPB VGND VPWR B1_N A2 X A1
X0 a_1021_47# A1 a_205_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X a_205_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 VPWR a_205_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_205_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND A2 a_1021_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND a_42_47# a_205_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_861_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.10075 ps=0.96 w=0.65 l=0.15
X7 a_205_21# A1 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.07475 ps=0.88 w=0.65 l=0.15
X8 X a_205_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_603_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND B1_N a_42_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.25025 ps=2.07 w=0.65 l=0.15
X11 VPWR A2 a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_603_297# a_42_47# a_205_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR a_205_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.15
X14 a_205_21# a_42_47# a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND a_205_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26325 pd=1.46 as=0.091 ps=0.93 w=0.65 l=0.15
X16 VPWR B1_N a_42_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X17 VGND a_205_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VPWR A1 a_603_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_603_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_205_21# a_42_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26325 ps=1.46 w=0.65 l=0.15
X21 X a_205_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND VNB VPB A_N B C D X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.10397 ps=1 w=0.65 l=0.15
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14325 pd=1.33 as=0.06615 ps=0.735 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10397 pd=1 as=0.06195 ps=0.715 w=0.42 l=0.15
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.09912 ps=0.955 w=0.65 l=0.15
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.14325 ps=1.33 w=1 l=0.15
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR VNB VPB X C B A_N
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12715 ps=1.095 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12715 pd=1.095 as=0.05355 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_4 VNB VPB VGND VPWR A2 A1 B1_N Y
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18362 ps=1.215 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18362 pd=1.215 as=0.16087 ps=1.145 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.16087 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 VPB VNB A1 A2 A3 Y B1 VPWR VGND
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 VNB VPB VGND VPWR Y B1 A2 A1 C1
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_2 VNB VPB VGND VPWR A2 A1 B1 B2 Y C1
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1755 ps=1.84 w=0.65 l=0.15
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 VPWR VGND VPB VNB A2 A1 Y B1 C1
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 VPB VNB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_4 VNB VPB VGND VPWR A_N X D C B
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_815_47# B a_701_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.1365 ps=1.07 w=0.65 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.135 ps=1.27 w=1 l=0.15
X5 a_174_21# a_27_47# a_815_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.143 ps=1.09 w=0.65 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_701_47# C a_617_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3275 ps=1.655 w=1 l=0.15
X10 a_174_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.21 ps=1.42 w=1 l=0.15
X11 VPWR a_27_47# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.22 ps=1.44 w=1 l=0.15
X12 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X13 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_617_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.21287 ps=1.305 w=0.65 l=0.15
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.21287 pd=1.305 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlxtn_2 VNB VPB VPWR VGND Q D GATE_N
X0 VPWR a_728_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_728_21# a_663_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2 VPWR a_728_21# a_686_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR GATE_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_686_413# a_27_47# a_565_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.09555 ps=0.875 w=0.42 l=0.15
X5 VGND a_728_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Q a_728_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X7 VGND a_565_413# a_728_21# VNB sky130_fd_pr__nfet_01v8 ad=0.09262 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_663_47# a_193_47# a_565_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0504 ps=0.64 w=0.36 l=0.15
X10 a_469_369# a_303_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0968 pd=0.97 as=0.0864 ps=0.91 w=0.64 l=0.15
X11 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 VPWR D a_303_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X14 a_565_413# a_193_47# a_469_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09555 pd=0.875 as=0.0968 ps=0.97 w=0.42 l=0.15
X15 VPWR a_565_413# a_728_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.26 ps=2.52 w=1 l=0.15
X16 a_469_47# a_303_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND GATE_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_565_413# a_27_47# a_469_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0504 pd=0.64 as=0.0777 ps=0.81 w=0.36 l=0.15
X19 Q a_728_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09262 ps=0.935 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s4s_1 VPWR VGND VPB VNB X A
X0 X a_345_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1 VPWR a_239_47# a_345_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND a_239_47# a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 X a_345_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 a_239_47# a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 a_239_47# a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR X a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND X a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_2 VNB VPB VGND VPWR A_N C B Y
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17575 pd=1.395 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11975 ps=1.045 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.17575 ps=1.395 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11975 pd=1.045 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VPB VGND VPWR VNB B1 X D1 A1 A2 C1
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.08287 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.27463 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.08287 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.27463 ps=1.495 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_4 VNB VPB VPWR VGND C1 Y B2 B1 A2 A1
X0 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X3 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X6 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X11 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.09425 pd=0.94 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X24 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X28 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09425 ps=0.94 w=0.65 l=0.15
X39 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt tt_um_femto VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7]
X_09671_ VGND VPWR VPWR VGND _14369_/D hold843/X _09687_/S fanout54/X sky130_fd_sc_hd__mux2_1
X_08622_ VGND VPWR VGND VPWR _15302_/D hold1079/X _08628_/A2 _08621_/X _11347_/A sky130_fd_sc_hd__o211a_1
X_08553_ VGND VPWR VGND VPWR _15315_/D hold1075/X _08553_/A2 _08552_/X _11431_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08484_ VPWR VGND VGND VPWR _08484_/X _15334_/Q _08484_/B sky130_fd_sc_hd__or2_1
X_07504_ VPWR VGND _07506_/A _07507_/B _15462_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_23_623 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07435_ VPWR VGND VGND VPWR _15457_/Q _07714_/A _07436_/B sky130_fd_sc_hd__nor2_1
X_12994__111 VPWR VGND VPWR VGND _14237_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
XFILLER_17_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07366_ VPWR VGND _08223_/B _07366_/B _07366_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_14105__1222 VPWR VGND VPWR VGND _15524_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_07297_ VPWR VGND VGND VPWR _15467_/Q _07297_/B _07860_/A sky130_fd_sc_hd__nor2_1
X_09105_ VGND VPWR VPWR VGND _14990_/D hold471/X _09124_/S clone55/X sky130_fd_sc_hd__mux2_1
X_09036_ VGND VPWR VPWR VGND _15054_/D hold346/X _09055_/S clone55/X sky130_fd_sc_hd__mux2_1
Xhold362 hold362/X hold362/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 hold351/X hold351/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 hold340/X hold340/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold373 hold373/X hold373/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold395 hold395/X hold395/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 hold384/X hold384/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ VPWR VGND VPWR VGND _14767_/Q _09938_/C _09938_/A _09939_/B sky130_fd_sc_hd__or3_1
Xfanout820 VPWR VGND _11308_/C1 fanout824/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout842 VGND VPWR _11341_/A _12751_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout831 VGND VPWR fanout844/X _12492_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout864 VGND VPWR _07119_/Y _07421_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout875 VGND VPWR _15582_/Q _08286_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout853 VPWR VGND _08240_/A _07966_/A VPWR VGND sky130_fd_sc_hd__buf_2
X_09869_ VPWR VGND VGND VPWR _09869_/A _09888_/S _09869_/B sky130_fd_sc_hd__nand2_1
Xhold1040 hold1040/X _14253_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout886 VPWR VGND _07141_/A _15573_/Q VPWR VGND sky130_fd_sc_hd__buf_2
Xhold1051 hold1051/X _14871_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13220__337 VPWR VGND VPWR VGND _14495_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_12880_ VPWR VGND VPWR VGND _08232_/Y _07574_/A _12878_/X _15603_/D sky130_fd_sc_hd__a21oi_1
X_11900_ VGND VPWR VGND VPWR _15453_/D _12195_/B1 _11898_/X _11899_/Y _11388_/S sky130_fd_sc_hd__o211a_1
Xhold1073 hold1073/X _14892_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 hold1084/X _14946_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 hold1062/X _14875_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ VPWR VGND VGND VPWR _11831_/X _12100_/S _11831_/B sky130_fd_sc_hd__or2_1
Xhold1095 hold1095/X _15021_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14550_ hold822/A _14550_/CLK _14550_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1298 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11762_ VGND VPWR VPWR VGND _11762_/X hold394/A _12086_/S hold240/A sky130_fd_sc_hd__mux2_1
X_14481_ hold912/A _14481_/CLK _14481_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11693_ VGND VPWR VPWR VGND _11693_/X _11690_/X _12476_/S _11689_/X sky130_fd_sc_hd__mux2_1
X_10713_ VGND VPWR VPWR VGND _10713_/X hold974/A _10743_/B hold422/A sky130_fd_sc_hd__mux2_1
X_13868__985 VPWR VGND VPWR VGND _15240_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
XFILLER_9_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10644_ VGND VPWR VPWR VGND _10644_/X _10641_/X _10652_/S _10640_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_148 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13114__231 VPWR VGND VPWR VGND _14357_/CLK clkload24/A sky130_fd_sc_hd__inv_2
XFILLER_31_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10575_ VGND VPWR VPWR VGND _10575_/X hold744/A _10730_/S hold444/A sky130_fd_sc_hd__mux2_1
X_15102_ _15102_/Q _15102_/CLK _15102_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12314_ VGND VPWR VPWR VGND _12314_/X _12311_/X _12684_/S _12310_/X sky130_fd_sc_hd__mux2_1
Xrebuffer7 VPWR VGND VPWR VGND _07477_/S rebuffer7/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15033_ hold653/A _15033_/CLK _15033_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12245_ VGND VPWR VPWR VGND _12245_/X hold493/A _12318_/S hold505/A sky130_fd_sc_hd__mux2_1
XFILLER_47_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12176_ VGND VPWR VPWR VGND _12177_/B _12175_/Y _12176_/S _12167_/Y sky130_fd_sc_hd__mux2_1
X_11127_ VGND VPWR VPWR VGND _11131_/B _14796_/Q _11146_/B _14247_/Q sky130_fd_sc_hd__mux2_1
XFILLER_7_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11058_ VGND VPWR VGND VPWR _11058_/X _11178_/C1 _11054_/X _11057_/X _11180_/C1 sky130_fd_sc_hd__o211a_1
X_10009_ VGND VPWR VPWR VGND _15619_/Q _15619_/D _10010_/C sky130_fd_sc_hd__xor2_1
XFILLER_75_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14817_ _14817_/Q clkload27/A _14817_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_64_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_910 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_75_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14748_ hold211/A _14748_/CLK _14748_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14679_ hold504/A _14679_/CLK _14679_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07220_ VGND VPWR VPWR VGND _07222_/A _07220_/S _15592_/Q _14381_/Q sky130_fd_sc_hd__mux2_4
X_07151_ VPWR VGND VGND VPWR _14409_/Q _07301_/A2 _07304_/B1 _07153_/B sky130_fd_sc_hd__o21a_1
X_07082_ VPWR VGND VPWR VGND _07082_/Y _07082_/A sky130_fd_sc_hd__inv_2
XFILLER_12_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13661__778 VPWR VGND VPWR VGND _15001_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_47_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout127 VGND VPWR _08190_/X _09827_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout105 VGND VPWR _09547_/A1 _08149_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout138 VPWR VGND _08700_/B1 _08730_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout116 VGND VPWR _09690_/A0 _08250_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout149 VGND VPWR _08686_/A2 _08613_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07984_ VGND VPWR VPWR VGND _07984_/X _10065_/C _07984_/S _12806_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09723_ VGND VPWR VPWR VGND _14320_/D _09723_/A1 _09728_/S hold689/X sky130_fd_sc_hd__mux2_1
X_09654_ VGND VPWR VPWR VGND _14416_/D hold816/X _09659_/S _09688_/A0 sky130_fd_sc_hd__mux2_1
X_08605_ VPWR VGND VGND VPWR _08605_/A _09001_/B _08605_/Y sky130_fd_sc_hd__nor2_1
Xtt_um_femto_898 uio_out[1] tt_um_femto_898/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09585_ VGND VPWR VPWR VGND _14480_/D hold864/X _09590_/S _09723_/A1 sky130_fd_sc_hd__mux2_1
X_13555__672 VPWR VGND VPWR VGND _14886_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_08536_ VPWR VGND VPWR VGND _08540_/B1 hold1414/X _08540_/A2 _08537_/B _15318_/Q
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08467_ VGND VPWR VGND VPWR _15343_/D hold1244/X _08483_/A2 _08466_/X _11974_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07418_ VPWR VGND VPWR VGND _07418_/B _08286_/B _10072_/A _07418_/X sky130_fd_sc_hd__or3_1
X_08398_ VGND VPWR VPWR VGND _15379_/D fanout21/X _08409_/S hold712/X sky130_fd_sc_hd__mux2_1
X_07349_ VGND VPWR VGND VPWR _07349_/X _07942_/B _07945_/A _07921_/A sky130_fd_sc_hd__a21bo_1
XFILLER_12_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10360_ VGND VPWR VPWR VGND _10360_/X hold919/A _10632_/B hold435/A sky130_fd_sc_hd__mux2_1
X_09019_ VPWR VGND VGND VPWR _09938_/A _09019_/B _15097_/D sky130_fd_sc_hd__nor2_1
X_10291_ VGND VPWR VPWR VGND _10291_/X hold778/A _10521_/B hold734/A sky130_fd_sc_hd__mux2_1
Xhold170 hold170/X hold170/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ VGND VPWR VPWR VGND _12030_/X hold887/A _12043_/B hold504/A sky130_fd_sc_hd__mux2_1
XFILLER_78_604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold181 hold181/X hold181/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/X hold192/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout650 VPWR VGND _09513_/S _09486_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout683 VPWR VGND _08375_/S _08366_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout672 _09194_/S _09164_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout694 VGND VPWR _08893_/A2 _08880_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout661 _09310_/S _09302_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12863_ VGND VPWR VPWR VGND _15587_/D _12863_/A1 _12870_/S hold1318/X sky130_fd_sc_hd__mux2_1
XFILLER_46_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14602_ _14602_/Q _14602_/CLK _14602_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11814_ VGND VPWR VGND VPWR _11814_/X _11813_/X _11812_/X _11810_/S _12748_/C1 sky130_fd_sc_hd__a211o_1
X_12794_ VPWR VGND VGND VPWR _12817_/A _12794_/Y _12794_/B sky130_fd_sc_hd__nand2_1
X_15582_ _15582_/Q clkload27/A _15582_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_26_280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14533_ hold157/A _14533_/CLK _14533_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11745_ VGND VPWR VGND VPWR _11745_/X _11742_/X _11744_/X _12720_/A1 _12415_/C1 sky130_fd_sc_hd__a211o_1
X_14464_ _14464_/Q _14464_/CLK _14464_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11676_ VPWR VGND _11676_/X _11675_/X _11671_/X _12176_/S _11667_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14395_ _14395_/Q clkload9/A _14395_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_31_1248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10627_ VGND VPWR VPWR VGND _10627_/X hold733/A _10627_/S hold300/A sky130_fd_sc_hd__mux2_1
X_10558_ VGND VPWR VGND VPWR _10558_/X _10662_/S _10553_/X _10557_/X _10667_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_6_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10489_ VPWR VGND VGND VPWR _10470_/Y _10488_/X _10192_/B _14389_/Q _14389_/D _08735_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12228_ VPWR VGND VGND VPWR _12228_/X hold622/A _12228_/B sky130_fd_sc_hd__or2_1
X_15016_ _15016_/Q _15016_/CLK _15016_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13498__615 VPWR VGND VPWR VGND _14773_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
XFILLER_2_880 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12159_ VPWR VGND VGND VPWR _12140_/Y _12158_/X _10562_/B _15460_/Q _15460_/D _12159_/C1
+ sky130_fd_sc_hd__o221a_1
X_14104__1221 VPWR VGND VPWR VGND _15523_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_13539__656 VPWR VGND VPWR VGND _14870_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_80_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09370_ VGND VPWR VPWR VGND _14676_/D hold836/X _09377_/S fanout7/X sky130_fd_sc_hd__mux2_1
X_08321_ VGND VPWR VPWR VGND _15498_/D fanout37/X _08330_/S hold926/X sky130_fd_sc_hd__mux2_1
X_08252_ VPWR VGND VPWR VGND _08174_/Y _15155_/Q _08252_/A2 _08252_/X _14837_/Q sky130_fd_sc_hd__a22o_1
XFILLER_60_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07203_ VPWR VGND VGND VPWR _08115_/A _07204_/B _08137_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08183_ VPWR VGND VPWR VGND _08293_/A3 _15071_/Q _08293_/B1 _08183_/X _07209_/X sky130_fd_sc_hd__a22o_1
X_07134_ VGND VPWR VPWR VGND _07765_/B _07807_/S _15574_/Q sky130_fd_sc_hd__and2b_2
XPHY_EDGE_ROW_58_Left_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_75_607 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07967_ VGND VPWR VGND VPWR _07983_/A _08007_/A _07982_/B _07981_/A sky130_fd_sc_hd__a21bo_1
X_09706_ VGND VPWR VPWR VGND _14337_/D _09710_/S fanout52/X hold1208/X sky130_fd_sc_hd__mux2_4
XFILLER_67_191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07898_ VPWR VGND VGND VPWR _07966_/A _07898_/Y _12822_/B sky130_fd_sc_hd__nand2_1
X_09637_ VGND VPWR VPWR VGND _14433_/D hold987/X _09637_/S clone5/A sky130_fd_sc_hd__mux2_1
X_13291__408 VPWR VGND VPWR VGND _14566_/CLK clkload53/A sky130_fd_sc_hd__inv_2
XFILLER_70_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09568_ VGND VPWR VPWR VGND _14497_/D _09584_/S hold1207/X clone46/X sky130_fd_sc_hd__mux2_4
XFILLER_3_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08519_ VPWR VGND VPWR VGND _08534_/B1 hold1460/X _08503_/A _08520_/B hold1416/X
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_67_Left_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09499_ VGND VPWR VPWR VGND _14560_/D _09517_/S fanout50/X hold1183/X sky130_fd_sc_hd__mux2_4
X_11530_ VGND VPWR VPWR VGND _11530_/X _11529_/X _11530_/S _15474_/Q sky130_fd_sc_hd__mux2_1
XFILLER_8_917 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13332__449 VPWR VGND VPWR VGND _14607_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_11461_ VGND VPWR VPWR VGND _11461_/X _11460_/X _11491_/S _15451_/Q sky130_fd_sc_hd__mux2_1
X_11392_ VPWR VGND VGND VPWR _14851_/Q _11393_/S _11392_/B sky130_fd_sc_hd__nand2_1
X_10412_ VGND VPWR VGND VPWR _10412_/X _10409_/X _10411_/X _10705_/A _10706_/C1 sky130_fd_sc_hd__a211o_1
X_14180_ hold642/A _14180_/CLK _14180_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10343_ VGND VPWR VPWR VGND _10343_/X hold969/A _10612_/S hold474/A sky130_fd_sc_hd__mux2_1
X_13185__302 VPWR VGND VPWR VGND _14460_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_76_Left_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10274_ VGND VPWR VPWR VGND _10274_/X _10271_/X _10613_/A _10270_/X sky130_fd_sc_hd__mux2_1
X_13226__343 VPWR VGND VPWR VGND _14501_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_12013_ VGND VPWR VPWR VGND _12013_/X hold763/A _12112_/S hold848/A sky130_fd_sc_hd__mux2_1
Xfanout491 VGND VPWR _11954_/S _11950_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout480 VGND VPWR _11628_/S _12089_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1293 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15634_ _15634_/Q clkload49/A _15634_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12846_ VPWR VGND _12846_/X _12846_/B _15571_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_15565_ _15565_/Q clkload50/A _15565_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_37_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12777_ VPWR VGND _12777_/X _12788_/S _08124_/X _08099_/B _12790_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_37_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14516_ hold158/A _14516_/CLK _14516_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11728_ VPWR VGND VGND VPWR _11728_/X _12396_/S _11728_/B sky130_fd_sc_hd__or2_1
X_15496_ hold936/A _15496_/CLK _15496_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11659_ VPWR VGND VGND VPWR _12029_/A _11659_/B _11659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_1192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14447_ hold693/A _14447_/CLK _14447_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14378_ _14378_/Q _14378_/CLK _14378_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold928 hold928/X hold928/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 hold917/X hold917/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold906 hold906/X hold906/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_3_1_0_clk clkload0/A clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold939 hold939/X hold939/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08870_ VPWR VGND VGND VPWR _08870_/X _15157_/Q _08918_/B sky130_fd_sc_hd__or2_1
X_07821_ VPWR VGND VGND VPWR _07857_/A _07821_/Y _10071_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07752_ VPWR VGND VPWR VGND _07751_/C _15597_/Q _15550_/Q _07753_/B sky130_fd_sc_hd__a21o_1
XFILLER_65_662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07683_ VPWR VGND VPWR VGND _07679_/Y _07328_/Y _07682_/X _07683_/Y sky130_fd_sc_hd__a21oi_1
X_09422_ VGND VPWR VPWR VGND _14630_/D _09443_/S clone47/X hold1195/X sky130_fd_sc_hd__mux2_4
XFILLER_53_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_80_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09353_ VGND VPWR VPWR VGND _14693_/D hold436/X _09357_/S fanout68/X sky130_fd_sc_hd__mux2_1
X_08304_ _09486_/B _08304_/X _09486_/A _09521_/A VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
X_09284_ VGND VPWR VPWR VGND _14757_/D fanout70/X _09304_/S hold296/X sky130_fd_sc_hd__mux2_1
X_08235_ VPWR VGND VPWR VGND _08174_/Y _15335_/Q _08253_/A2 _08235_/X _14838_/Q sky130_fd_sc_hd__a22o_1
XFILLER_60_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13667__784 VPWR VGND VPWR VGND _15007_/CLK clkload19/A sky130_fd_sc_hd__inv_2
X_08166_ VPWR VGND VPWR VGND _08162_/A _08280_/A2 _08166_/X _08293_/B1 _15072_/Q _08165_/X
+ sky130_fd_sc_hd__a221o_1
X_07117_ VPWR VGND VPWR VGND _07827_/C _12878_/A sky130_fd_sc_hd__inv_2
XFILLER_10_1129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08097_ VGND VPWR _08097_/B _12781_/A _08097_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_12954__71 VPWR VGND VPWR VGND _14197_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
XFILLER_69_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08999_ VGND VPWR VGND VPWR _08999_/X _09007_/A _08937_/Y _15103_/Q _08998_/Y sky130_fd_sc_hd__a211o_1
XFILLER_21_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10961_ VPWR VGND VGND VPWR _10961_/X hold156/A _11142_/S sky130_fd_sc_hd__or2_1
X_12700_ VGND VPWR VGND VPWR _12700_/X hold932/A _12705_/A2 _12256_/S _12699_/X sky130_fd_sc_hd__o211a_1
X_10892_ VPWR VGND VGND VPWR _10889_/X _10891_/X _10987_/S _10892_/X sky130_fd_sc_hd__o21a_1
X_12631_ VPWR VGND VGND VPWR _12631_/X hold263/A _12736_/B sky130_fd_sc_hd__or2_1
XFILLER_19_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15350_ _15350_/Q _15350_/CLK _15350_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12562_ VGND VPWR VPWR VGND _12562_/X hold698/A _12671_/S hold306/A sky130_fd_sc_hd__mux2_1
X_14301_ hold183/A _14301_/CLK _14301_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11513_ VGND VPWR VPWR VGND _15088_/D _11512_/X _11538_/S _15088_/Q sky130_fd_sc_hd__mux2_1
X_15281_ _15281_/Q _15281_/CLK _15281_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12493_ VGND VPWR VPWR VGND _12497_/B hold579/A _12664_/S hold592/A sky130_fd_sc_hd__mux2_1
X_11444_ VGND VPWR VPWR VGND _15065_/D _11443_/Y _11477_/S hold1317/X sky130_fd_sc_hd__mux2_1
X_14232_ hold302/A _14232_/CLK _14232_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14103__1220 VPWR VGND VPWR VGND _15522_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_14193__911 _14193_/D _14193__911/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_14163_ hold506/A _14163_/CLK _14163_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11375_ VGND VPWR VPWR VGND _11375_/X _11374_/X _11387_/S _14846_/Q sky130_fd_sc_hd__mux2_1
X_10326_ VGND VPWR VPWR VGND _10326_/X _14868_/Q _11261_/B hold315/A sky130_fd_sc_hd__mux2_1
X_10257_ VGND VPWR VPWR VGND _10257_/X hold755/A _10258_/B hold511/A sky130_fd_sc_hd__mux2_1
X_13460__577 VPWR VGND VPWR VGND _14735_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_10188_ VGND VPWR VGND VPWR _10188_/X _10703_/A _10184_/X _10187_/X _10706_/C1 sky130_fd_sc_hd__o211a_1
X_14996_ hold340/A _14996_/CLK _14996_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15617_ _15617_/Q clkload27/A _15617_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12829_ VGND VPWR VPWR VGND _12830_/B _07865_/B _12829_/S _07869_/B sky130_fd_sc_hd__mux2_1
X_15548_ _15548_/Q clkload43/A _15548_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13354__471 VPWR VGND VPWR VGND _14629_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_15479_ _15479_/Q _15479_/CLK _15479_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08020_ VGND VPWR _07998_/C _08019_/X _08020_/Y _07733_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_50_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold703 hold703/X hold703/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold714 hold714/X hold714/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 hold725/X hold725/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 hold736/X hold736/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout7 VPWR VGND fanout7/X fanout7/A VPWR VGND sky130_fd_sc_hd__buf_6
X_09971_ VPWR VGND _15480_/D _09970_/Y _09890_/A _09977_/A _09969_/X VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold769 hold769/X hold769/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 hold758/X hold758/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13701__818 VPWR VGND VPWR VGND _15041_/CLK clkload22/A sky130_fd_sc_hd__inv_2
Xhold747 hold747/X hold747/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ VPWR VGND VGND VPWR _08922_/X _08922_/A _08924_/B sky130_fd_sc_hd__or2_1
Xhold1425 hold1425/X _15125_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 hold1414/X _15317_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08853_ VPWR VGND VGND VPWR _08853_/A _08853_/B _08853_/Y sky130_fd_sc_hd__nor2_1
Xhold1403 _09977_/B _14801_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 hold1447/X _15125_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 hold1436/X _15320_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07804_ VGND VPWR VGND VPWR _07888_/B _07909_/A _07803_/B _07803_/A sky130_fd_sc_hd__a21bo_1
Xhold1458 hold1458/X _15628_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08784_ VGND VPWR VPWR VGND _15225_/D fanout85/X _08808_/S hold222/X sky130_fd_sc_hd__mux2_1
Xhold1469 _08922_/A _15131_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07735_ VPWR VGND VPWR VGND _07827_/D _08286_/A _07714_/X _07736_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07666_ VPWR VGND VGND VPWR _07652_/B _07665_/Y _07984_/S _07666_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09405_ VGND VPWR VPWR VGND _14644_/D hold481/X _09406_/S fanout6/X sky130_fd_sc_hd__mux2_1
X_07597_ VGND VPWR VGND VPWR _07597_/X _10072_/A _07596_/X _07570_/X _07574_/A sky130_fd_sc_hd__o211a_4
XFILLER_0_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09336_ VGND VPWR VPWR VGND _14708_/D hold674/X _09336_/S fanout7/X sky130_fd_sc_hd__mux2_1
X_09267_ VGND VPWR VPWR VGND _14776_/D _09825_/A1 _09275_/S hold811/X sky130_fd_sc_hd__mux2_1
X_08218_ VGND VPWR _08218_/B _08218_/Y _08218_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_09198_ VGND VPWR VGND VPWR _09198_/X _09164_/A _09198_/C _09198_/B _15577_/Q sky130_fd_sc_hd__or4b_4
X_08149_ VGND VPWR VGND VPWR _08149_/X _08134_/Y _07996_/X _08143_/X _08148_/X sky130_fd_sc_hd__a211o_2
X_11160_ VPWR VGND VGND VPWR _11160_/X _11170_/S _11160_/B sky130_fd_sc_hd__or2_1
X_14218__936 _14218_/D _14218__936/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_11091_ VGND VPWR VPWR VGND _11091_/X _14470_/Q _11091_/S _14758_/Q sky130_fd_sc_hd__mux2_1
XFILLER_27_1412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10111_ VGND VPWR VGND VPWR _10111_/X hold956/A _10629_/A2 _10110_/X _10510_/S sky130_fd_sc_hd__o211a_1
X_10042_ VPWR VGND VGND VPWR _10042_/A _10042_/B _10043_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_49_927 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14850_ _14850_/Q clkload19/A _14850_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13297__414 VPWR VGND VPWR VGND _14572_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_14781_ hold574/A _14781_/CLK _14781_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11993_ VGND VPWR VPWR VGND _11993_/X _14422_/Q _11998_/S hold815/A sky130_fd_sc_hd__mux2_1
X_13338__455 VPWR VGND VPWR VGND _14613_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_10944_ VGND VPWR VPWR VGND _10944_/X _14210_/Q _11167_/S hold174/A sky130_fd_sc_hd__mux2_1
X_10875_ VGND VPWR VGND VPWR _10875_/X _12868_/A1 _10870_/X _10874_/X _10987_/S sky130_fd_sc_hd__o211a_1
XFILLER_34_1405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12614_ VGND VPWR VPWR VGND _12614_/X _14215_/Q _12635_/B _15223_/Q sky130_fd_sc_hd__mux2_1
X_15402_ hold556/A _15402_/CLK _15402_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15333_ _15333_/Q _15333_/CLK _15333_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12545_ VPWR VGND VPWR VGND _12544_/X _12656_/A1 _12543_/X _12545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15264_ _15264_/Q _15264_/CLK _15264_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12476_ VGND VPWR VPWR VGND _12476_/X _12475_/X _12476_/S _12474_/X sky130_fd_sc_hd__mux2_1
X_11427_ VGND VPWR VGND VPWR _14928_/D _14929_/Q _11431_/A2 _11426_/X _11431_/C1 sky130_fd_sc_hd__o211a_1
XANTENNA_5 _07631_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_15195_ hold224/A _15195_/CLK _15195_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14215_ _14215_/Q _14215_/CLK _14215_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14146_ _14146_/Q _14146_/CLK _14146_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11358_ VGND VPWR VPWR VGND _14857_/Q _14859_/Q _14858_/Q _11359_/C sky130_fd_sc_hd__or3b_1
X_10309_ VGND VPWR VGND VPWR _10309_/X hold805/A _11262_/A2 _10308_/X _11112_/A sky130_fd_sc_hd__o211a_1
XFILLER_80_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11289_ VGND VPWR VPWR VGND _11290_/B _14813_/Q _11299_/S _14381_/Q sky130_fd_sc_hd__mux2_1
XFILLER_67_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_67_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07520_ VPWR VGND VPWR VGND _07518_/X _07429_/A _07519_/Y _07526_/A sky130_fd_sc_hd__a21oi_1
Xrebuffer39 VPWR VGND VPWR VGND rebuffer39/X rebuffer40/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer28 VPWR VGND VPWR VGND rebuffer28/X rebuffer29/X sky130_fd_sc_hd__dlygate4sd1_1
X_14979_ hold899/A _14979_/CLK _14979_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_643 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07451_ VPWR VGND VPWR VGND _08580_/A _07452_/B sky130_fd_sc_hd__inv_2
XFILLER_50_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_22_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07382_ VPWR VGND VPWR VGND _07379_/X _07088_/Y _07258_/B _08026_/B _07381_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13090__207 VPWR VGND VPWR VGND _14333_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_09121_ VGND VPWR VPWR VGND _14974_/D hold524/X _09128_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_09052_ VGND VPWR VPWR VGND _15038_/D hold747/X _09059_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_13131__248 VPWR VGND VPWR VGND _14374_/CLK clkload48/A sky130_fd_sc_hd__inv_2
Xhold500 hold500/X hold500/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08003_ VGND VPWR _07272_/C _07272_/D _08025_/B _08041_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold511 hold511/X hold511/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 hold522/X hold522/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 hold533/X hold533/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 hold544/X hold544/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 hold588/X hold588/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 hold577/X hold577/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12924__41 VPWR VGND VPWR VGND _14167_/CLK clkload9/A sky130_fd_sc_hd__inv_2
Xhold566 hold566/X hold566/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 hold555/X hold555/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ VPWR VGND VPWR VGND _09954_/B _09954_/C _14127_/Q _09954_/X sky130_fd_sc_hd__or3_1
Xhold599 hold599/X hold599/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09885_ VPWR VGND VPWR VGND _14148_/Q _09885_/C hold212/A _09886_/B sky130_fd_sc_hd__or3_1
X_08905_ VGND VPWR VGND VPWR _15140_/D hold1373/X _08880_/B _08904_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
X_13779__896 VPWR VGND VPWR VGND _15151_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
Xhold1200 hold1200/X _14881_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 hold1233/X _15338_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 _14835_/D _11348_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1222 hold1222/X _14368_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ VGND VPWR VPWR VGND _15177_/D fanout25/X _08850_/S hold407/X sky130_fd_sc_hd__mux2_1
Xhold1255 hold1255/X _14841_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 hold1266/X _14470_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 hold1244/X _15342_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13025__142 VPWR VGND VPWR VGND _14268_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
Xhold1288 hold1288/X _15440_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 hold1277/X _15135_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 hold1299/X _14849_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ VGND VPWR VPWR VGND _15239_/D fanout15/X _08779_/S hold187/X sky130_fd_sc_hd__mux2_1
X_07718_ VPWR VGND VGND VPWR _07718_/A _07718_/B _07915_/A sky130_fd_sc_hd__nor2_1
X_08698_ VGND VPWR VGND VPWR _15282_/D hold978/X _08701_/A2 _08697_/X _12233_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_53_462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07649_ VPWR VGND VGND VPWR _07664_/A _07653_/A _07668_/A _07649_/Y sky130_fd_sc_hd__nor3_1
X_10660_ VGND VPWR VPWR VGND _10660_/X hold874/A _10720_/S hold558/A sky130_fd_sc_hd__mux2_1
XFILLER_41_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09319_ VGND VPWR VPWR VGND _14725_/D hold708/X _09327_/S fanout69/X sky130_fd_sc_hd__mux2_1
X_10591_ VPWR VGND VGND VPWR _10591_/X hold155/A _10742_/S sky130_fd_sc_hd__or2_1
X_12330_ VGND VPWR VGND VPWR _12330_/X hold817/A _12705_/A2 _12588_/A1 _12329_/X sky130_fd_sc_hd__o211a_1
X_12261_ VGND VPWR VPWR VGND _12261_/X hold770/A _12339_/B hold311/A sky130_fd_sc_hd__mux2_1
X_13723__840 VPWR VGND VPWR VGND _15063_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_11212_ VGND VPWR VPWR VGND _11212_/X hold980/A _11216_/S hold911/A sky130_fd_sc_hd__mux2_1
X_12192_ VGND VPWR VGND VPWR _12192_/X _15015_/Q _12192_/A2 _12180_/S _12191_/X sky130_fd_sc_hd__o211a_1
X_11143_ VGND VPWR VPWR VGND _11143_/X _11142_/X _11143_/S _11141_/X sky130_fd_sc_hd__mux2_1
X_11074_ VGND VPWR VGND VPWR _11074_/X _11071_/X _11073_/X _11185_/A1 _11254_/C1 sky130_fd_sc_hd__a211o_1
X_10025_ VPWR VGND VPWR VGND _10024_/C _15625_/Q hold1333/X _10025_/Y sky130_fd_sc_hd__a21oi_1
X_14902_ hold344/A _14902_/CLK _14902_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_223 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_267 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14833_ _14833_/Q clkload30/A _14833_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14764_ hold148/A _14764_/CLK _14764_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11976_ VGND VPWR VPWR VGND _11976_/X hold795/A _12006_/B hold651/A sky130_fd_sc_hd__mux2_1
XFILLER_44_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13572__689 VPWR VGND VPWR VGND _14903_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_14695_ hold487/A _14695_/CLK _14695_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10927_ VGND VPWR VPWR VGND _10927_/X hold428/A _11240_/S hold688/A sky130_fd_sc_hd__mux2_1
X_10858_ VPWR VGND VGND VPWR _10858_/X _14399_/Q _12269_/B sky130_fd_sc_hd__or2_1
X_10789_ VPWR VGND VGND VPWR _10789_/X hold321/A _11204_/S sky130_fd_sc_hd__or2_1
X_15316_ _15316_/Q _15316_/CLK _15316_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12528_ VPWR VGND VPWR VGND _12527_/X _12658_/A _12750_/B1 _12528_/X sky130_fd_sc_hd__a21o_1
X_15247_ hold317/A _15247_/CLK _15247_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12459_ VGND VPWR VPWR VGND _12459_/X hold516/A _12477_/B hold269/A sky130_fd_sc_hd__mux2_1
X_13466__583 VPWR VGND VPWR VGND _14741_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_15178_ hold393/A _15178_/CLK _15178_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14129_ _14129_/Q _14129_/CLK _14129_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout309 VPWR VGND _10553_/S fanout314/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_80_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13009__126 VPWR VGND VPWR VGND _14252_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_09670_ VGND VPWR VPWR VGND _14370_/D hold866/X _09687_/S clone54/X sky130_fd_sc_hd__mux2_1
X_08621_ VGND VPWR VGND VPWR _08621_/X _08626_/A _08627_/C1 hold940/X _08620_/Y sky130_fd_sc_hd__a211o_1
XFILLER_55_749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08552_ VGND VPWR VGND VPWR _08552_/X _08562_/A _08615_/B1 hold942/A _08551_/Y sky130_fd_sc_hd__a211o_1
XFILLER_78_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08483_ VGND VPWR VGND VPWR _15335_/D hold1286/X _08483_/A2 _08482_/X _11431_/C1
+ sky130_fd_sc_hd__o211a_1
X_07503_ VPWR VGND VGND VPWR _07531_/C _07530_/C _07503_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_996 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_35_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_23_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07434_ VPWR VGND _08544_/A _15601_/Q _15457_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_17_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07365_ VGND VPWR VGND VPWR _07366_/B _08275_/A _10061_/A _08258_/B _10062_/A sky130_fd_sc_hd__a211o_1
X_07296_ VPWR VGND VPWR VGND _07296_/Y _07298_/A sky130_fd_sc_hd__inv_2
X_09104_ VGND VPWR VPWR VGND _14991_/D hold301/X _09125_/S fanout63/X sky130_fd_sc_hd__mux2_1
X_13707__824 VPWR VGND VPWR VGND _15047_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_09035_ VGND VPWR VPWR VGND _15055_/D hold542/X _09056_/S fanout63/X sky130_fd_sc_hd__mux2_1
Xhold352 hold352/X hold352/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 hold341/X hold341/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 hold330/X hold330/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 hold374/X hold374/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 hold385/X hold385/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 hold396/X hold396/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 hold363/X hold363/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout821 VPWR VGND _08541_/A fanout824/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout810 VGND VPWR _08735_/C _08529_/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout832 VPWR VGND _11327_/A _09000_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout843 VPWR VGND _11341_/A fanout844/X VPWR VGND sky130_fd_sc_hd__buf_4
X_09937_ VPWR VGND VGND VPWR _09937_/A _09937_/B _14763_/D _09937_/Y sky130_fd_sc_hd__nor3_2
Xfanout876 VPWR VGND _09240_/A _15581_/Q VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout865 VPWR VGND _07418_/B _07119_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout854 VGND VPWR _07328_/Y _07966_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09868_ _09869_/B _09890_/A _15479_/Q _15477_/Q _09977_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xfanout887 VGND VPWR _10056_/A _10060_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold1041 hold1041/X _14874_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1030 hold1030/X _14484_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _11539_/B _14800_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 hold1052/X _15306_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 hold1063/X _15305_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ VPWR VGND VGND VPWR _09799_/B _09799_/Y _09799_/A sky130_fd_sc_hd__nor2_2
X_08819_ _15194_/D fanout93/X fanout89/X _08817_/Y _08818_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_2_1222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1074 hold1074/X _14890_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ VGND VPWR VPWR VGND _11830_/X hold665/A _12171_/S hold173/A sky130_fd_sc_hd__mux2_1
Xhold1096 hold1096/X _14664_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11761_ VGND VPWR VPWR VGND _11765_/B hold534/A _12086_/S hold229/A sky130_fd_sc_hd__mux2_1
X_10712_ VGND VPWR VPWR VGND _10716_/B hold618/A _10743_/B hold319/A sky130_fd_sc_hd__mux2_1
XFILLER_70_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11692_ VGND VPWR VGND VPWR _11692_/X _12489_/A1 _11688_/X _11691_/X _12485_/C1 sky130_fd_sc_hd__o211a_1
X_14480_ hold864/A _14480_/CLK _14480_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10643_ VGND VPWR VGND VPWR _10643_/X _10557_/A _10639_/X _10642_/X _10717_/C1 sky130_fd_sc_hd__o211a_1
X_10574_ VGND VPWR VPWR VGND _10574_/X _14200_/Q _10730_/S hold181/A sky130_fd_sc_hd__mux2_1
X_13153__270 VPWR VGND VPWR VGND _14428_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_15101_ hold971/A _15101_/CLK hold972/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12313_ VGND VPWR VGND VPWR _12313_/X _12580_/A1 _12309_/X _12312_/X _12702_/C1 sky130_fd_sc_hd__o211a_1
Xrebuffer8 VPWR VGND VPWR VGND _07826_/A _07477_/S sky130_fd_sc_hd__dlygate4sd1_1
X_15032_ hold727/A _15032_/CLK _15032_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12244_ VGND VPWR VPWR VGND _12244_/X _12243_/X _12581_/S _12242_/X sky130_fd_sc_hd__mux2_1
X_12175_ VPWR VGND VPWR VGND _12174_/X _12175_/A1 _12173_/X _12175_/Y sky130_fd_sc_hd__a21oi_1
X_11126_ VPWR VGND VPWR VGND _11125_/X _11245_/A1 _11124_/X _11126_/Y sky130_fd_sc_hd__a21oi_1
X_13500__617 VPWR VGND VPWR VGND _14775_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
XFILLER_49_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11057_ VPWR VGND VGND VPWR _11057_/X _11176_/S _11057_/B sky130_fd_sc_hd__or2_1
XFILLER_7_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10008_ VPWR VGND VGND VPWR _10010_/C _10008_/B _15618_/D sky130_fd_sc_hd__nor2_1
X_14816_ _14816_/Q clkload20/A _14816_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11959_ VGND VPWR VGND VPWR _11959_/X _11948_/S _11954_/X _11958_/X _12189_/C1 sky130_fd_sc_hd__o211a_1
X_14747_ hold242/A _14747_/CLK _14747_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_33_933 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_60_774 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14678_ hold815/A _14678_/CLK _14678_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1190 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07150_ VPWR VGND VGND VPWR _07411_/A _07416_/A _08287_/A sky130_fd_sc_hd__nor2_2
XFILLER_12_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout106 VGND VPWR _12829_/S _12788_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout128 VPWR VGND _09826_/A1 _09548_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout117 VGND VPWR _09655_/A0 _09863_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09722_ VGND VPWR VPWR VGND _14321_/D _09827_/A1 _09725_/S hold805/X sky130_fd_sc_hd__mux2_1
X_07983_ VPWR VGND VGND VPWR _07983_/A _10065_/C _07983_/B sky130_fd_sc_hd__nand2_1
Xfanout139 VGND VPWR _08730_/B1 _08688_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_55_535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09653_ VGND VPWR VPWR VGND _14417_/D hold962/X _09656_/S _09653_/A0 sky130_fd_sc_hd__mux2_1
X_09584_ VGND VPWR VPWR VGND _14481_/D hold912/X _09584_/S _09827_/A1 sky130_fd_sc_hd__mux2_1
X_08604_ VGND VPWR VPWR VGND _09001_/B _15549_/Q _07552_/B1 _08604_/B2 _08603_/Y sky130_fd_sc_hd__o2bb2a_1
Xtt_um_femto_899 uio_out[2] tt_um_femto_899/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08535_ VPWR VGND _15319_/D _08535_/B _08541_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_13096__213 VPWR VGND VPWR VGND _14339_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_08466_ VPWR VGND VGND VPWR _08466_/X _08466_/A _08482_/B sky130_fd_sc_hd__or2_1
XFILLER_51_763 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07417_ _08286_/B _08286_/A _07417_/X _15584_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_08397_ VGND VPWR VPWR VGND _15380_/D fanout26/X _08411_/S hold733/X sky130_fd_sc_hd__mux2_1
X_14062__1179 VPWR VGND VPWR VGND _15481_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_13137__254 VPWR VGND VPWR VGND _14412_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_07348_ VPWR VGND VGND VPWR _07285_/B _15463_/Q _07921_/A sky130_fd_sc_hd__nand2b_1
XFILLER_12_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07279_ VPWR VGND VPWR VGND _07279_/Y _07926_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09018_ VPWR VGND VPWR VGND _08937_/Y hold928/X _08933_/A _09019_/B sky130_fd_sc_hd__a21oi_1
XFILLER_3_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10290_ VGND VPWR VGND VPWR _10290_/X hold856/A _10633_/A2 _10289_/X _10523_/A1 sky130_fd_sc_hd__o211a_1
Xhold160 hold160/X hold160/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold171/X hold171/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold182/X hold182/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13794__911 VPWR VGND VPWR VGND _15166_/CLK clkload37/A sky130_fd_sc_hd__inv_2
Xhold193 hold193/X hold193/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout651 _09514_/S _09517_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_59_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout640 _09590_/S _09588_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout673 _09128_/S _09126_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_24_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout662 VPWR VGND _09302_/S _09276_/Y VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_8_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout684 VPWR VGND _08366_/S _08342_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout695 VPWR VGND _08893_/A2 _08863_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_13835__952 VPWR VGND VPWR VGND _15207_/CLK clkload20/A sky130_fd_sc_hd__inv_2
XFILLER_19_738 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12862_ VGND VPWR VPWR VGND _15586_/D _12367_/S _12870_/S hold1329/X sky130_fd_sc_hd__mux2_1
X_11813_ VGND VPWR VPWR VGND _11813_/X _14868_/Q _12747_/S hold315/A sky130_fd_sc_hd__mux2_1
X_14601_ hold234/A _14601_/CLK _14601_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15581_ _15581_/Q clkload31/A _15581_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12793_ VPWR VGND _12793_/X _12820_/B _08038_/X _07837_/Y _12792_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_42_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14532_ hold295/A _14532_/CLK _14532_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11744_ VGND VPWR VGND VPWR _11744_/X _15003_/Q _12488_/A2 _12721_/S _11743_/X sky130_fd_sc_hd__o211a_1
X_14463_ hold573/A _14463_/CLK _14463_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11675_ VGND VPWR VGND VPWR _11675_/X _11672_/X _11674_/X _11894_/S _12185_/A1 sky130_fd_sc_hd__a211o_1
X_10626_ VGND VPWR VGND VPWR _10626_/X _10634_/C1 _10625_/X _10622_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
X_14394_ _14394_/Q clkload18/A _14394_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10557_ VPWR VGND VGND VPWR _10557_/X _10557_/A _10557_/B sky130_fd_sc_hd__or2_1
X_10488_ VPWR VGND VPWR VGND _10487_/X _10507_/A _12195_/B1 _10488_/X sky130_fd_sc_hd__a21o_1
X_15015_ _15015_/Q _15015_/CLK _15015_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12227_ VGND VPWR VPWR VGND _12227_/X hold646/A _12227_/S hold595/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12158_ VPWR VGND VPWR VGND _12157_/X _12214_/A _11973_/B _12158_/X sky130_fd_sc_hd__a21o_1
X_11109_ VGND VPWR VPWR VGND _11109_/X _15393_/Q _11109_/S _15540_/Q sky130_fd_sc_hd__mux2_1
X_12089_ VGND VPWR VPWR VGND _12089_/X _14553_/Q _12089_/S hold245/A sky130_fd_sc_hd__mux2_1
X_13578__695 VPWR VGND VPWR VGND _14909_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_42_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08320_ VGND VPWR VPWR VGND _15499_/D fanout38/X _08332_/S hold770/X sky130_fd_sc_hd__mux2_1
XFILLER_33_752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08251_ VGND VPWR VPWR VGND _15516_/D _09228_/A0 _08251_/S hold290/X sky130_fd_sc_hd__mux2_1
X_07202_ VPWR VGND VGND VPWR _15453_/Q _07358_/B _07204_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15266__941 _15266_/D _15266__941/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08182_ VGND VPWR VPWR VGND _08182_/X _08181_/X _08182_/S _12766_/B sky130_fd_sc_hd__mux2_1
X_07133_ VPWR VGND VPWR VGND _07133_/Y _08231_/S sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_1256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13819__936 VPWR VGND VPWR VGND _15191_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_07966_ VPWR VGND VGND VPWR _07966_/A _07966_/Y _12810_/B sky130_fd_sc_hd__nand2_1
X_09705_ VGND VPWR VPWR VGND _14338_/D fanout57/X _09710_/S hold713/X sky130_fd_sc_hd__mux2_1
X_07897_ VPWR VGND VGND VPWR _07897_/A _12822_/B _07897_/B sky130_fd_sc_hd__nand2_1
X_09636_ VGND VPWR VPWR VGND _14434_/D hold774/X _09637_/S clone54/X sky130_fd_sc_hd__mux2_1
XFILLER_56_899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_43_505 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09567_ VGND VPWR VPWR VGND _14498_/D hold787/X _09584_/S clone54/X sky130_fd_sc_hd__mux2_1
X_08518_ VPWR VGND _15327_/D _08518_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
X_09498_ VGND VPWR VPWR VGND _14561_/D _09514_/S fanout52/X hold1270/X sky130_fd_sc_hd__mux2_4
X_08449_ VGND VPWR VGND VPWR _15352_/D hold1327/X _08448_/B _08448_/Y _11399_/A1 sky130_fd_sc_hd__o211a_1
X_13371__488 VPWR VGND VPWR VGND _14646_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_11460_ VGND VPWR VPWR VGND _11460_/X _15072_/Q _11475_/S _15070_/Q sky130_fd_sc_hd__mux2_1
XFILLER_17_1082 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11391_ VPWR VGND VPWR VGND _11387_/S _09938_/A hold1335/X _14850_/D _11390_/X sky130_fd_sc_hd__a22o_1
X_10411_ VGND VPWR VGND VPWR _10411_/X _15007_/Q _10688_/A2 _10410_/X _10703_/A sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10342_ VGND VPWR VPWR VGND _10346_/B hold462/A _10353_/S hold350/A sky130_fd_sc_hd__mux2_1
X_12012_ VGND VPWR VPWR VGND _12016_/B hold547/A _12112_/S hold472/A sky130_fd_sc_hd__mux2_1
X_10273_ VGND VPWR VGND VPWR _10273_/X _10614_/A1 _10269_/X _10272_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
X_13265__382 VPWR VGND VPWR VGND _14540_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_8_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout492 VGND VPWR _11954_/S _11964_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_65_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout470 VGND VPWR _12080_/A2 _12743_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout481 VGND VPWR fanout497/X _11628_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_15702_ VGND VPWR _15702_/A uo_out[7] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_46_343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_1158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15633_ _15633_/Q clkload49/A _15633_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12845_ VPWR VGND _12845_/X _12845_/B _12845_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_62_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15564_ _15564_/Q clkload44/A _15564_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12776_ VPWR VGND VGND VPWR _12776_/A _12788_/S _12776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13612__729 VPWR VGND VPWR VGND _14952_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_14515_ hold381/A _14515_/CLK _14515_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11727_ VGND VPWR VPWR VGND _11727_/X hold693/A _11748_/S hold281/A sky130_fd_sc_hd__mux2_1
X_15495_ hold917/A _15495_/CLK _15495_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11658_ VGND VPWR VPWR VGND _11659_/B _11657_/Y _12176_/S _11649_/Y sky130_fd_sc_hd__mux2_1
X_14446_ hold937/A _14446_/CLK _14446_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14377_ hold980/A _14377_/CLK _14377_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11589_ VPWR VGND VGND VPWR _11589_/X hold369/A _11756_/S sky130_fd_sc_hd__or2_1
X_10609_ VGND VPWR VPWR VGND _10613_/B hold384/A _10609_/S hold184/A sky130_fd_sc_hd__mux2_1
Xhold907 hold907/X hold907/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 hold918/X hold918/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 hold929/X hold929/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13506__623 VPWR VGND VPWR VGND _14781_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
XFILLER_43_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14061__1178 VPWR VGND VPWR VGND _15480_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_07820_ VGND VPWR _10071_/B _07820_/A _07820_/B VPWR VGND sky130_fd_sc_hd__xnor2_2
X_07751_ VGND VPWR _07751_/X _15597_/Q _15550_/Q _07751_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_65_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07682_ VPWR VGND VPWR VGND _07681_/Y _07857_/A _07333_/Y _07682_/X sky130_fd_sc_hd__a21o_1
X_09421_ VGND VPWR VPWR VGND _14631_/D fanout78/X _09443_/S hold629/X sky130_fd_sc_hd__mux2_1
XFILLER_80_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09352_ VGND VPWR VPWR VGND _14694_/D hold570/X _09357_/S _07659_/X sky130_fd_sc_hd__mux2_1
X_08303_ VPWR VGND _09557_/A _09486_/B _09164_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_09283_ VGND VPWR VPWR VGND _14758_/D _09304_/S fanout74/X hold1155/X sky130_fd_sc_hd__mux2_4
X_08234_ VPWR VGND VGND VPWR _07645_/X _08232_/Y _08072_/X _08233_/X _08234_/X sky130_fd_sc_hd__o22a_1
X_08165_ VPWR VGND VGND VPWR _15452_/Q _07371_/B _08278_/B _08165_/X sky130_fd_sc_hd__o21a_1
X_07116_ VPWR VGND VPWR VGND _07827_/B _15572_/Q sky130_fd_sc_hd__inv_2
X_08096_ VPWR VGND VGND VPWR _08096_/A _08096_/B _08097_/B sky130_fd_sc_hd__nor2_1
X_13249__366 VPWR VGND VPWR VGND _14524_/CLK clkload17/A sky130_fd_sc_hd__inv_2
XFILLER_76_939 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08998_ VPWR VGND VGND VPWR _09007_/A _08998_/B _08998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07949_ VGND VPWR _07962_/A _07950_/A _15561_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_67_clk _12955__72/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_29_877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10960_ VGND VPWR VPWR VGND _10960_/X hold687/A _11142_/S hold162/A sky130_fd_sc_hd__mux2_1
XFILLER_71_644 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10891_ VGND VPWR VGND VPWR _10891_/X _10333_/A _10886_/X _10890_/X _10891_/C1 sky130_fd_sc_hd__o211a_1
X_09619_ VGND VPWR VPWR VGND _14449_/D _09653_/A0 _09619_/S hold862/X sky130_fd_sc_hd__mux2_1
X_12630_ VGND VPWR VPWR VGND _12630_/X hold537/A _12736_/B hold655/A sky130_fd_sc_hd__mux2_1
XFILLER_58_1182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12561_ VGND VPWR VGND VPWR _12561_/X _15507_/Q _12669_/A2 _12735_/S _12560_/X sky130_fd_sc_hd__o211a_1
XFILLER_11_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11512_ VGND VPWR VPWR VGND _11512_/X _11511_/X _11530_/S _15468_/Q sky130_fd_sc_hd__mux2_1
X_15280_ _15280_/Q _15280_/CLK _15280_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14300_ hold408/A _14300_/CLK _14300_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12492_ VPWR VGND VGND VPWR _12473_/Y _12491_/X _12380_/B _15469_/Q _15469_/D _12492_/C1
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14231_ hold175/A _14231_/CLK _14231_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11443_ VPWR VGND VPWR VGND _12845_/B _08290_/A _11442_/Y _11443_/Y sky130_fd_sc_hd__a21oi_1
X_14162_ hold474/A _14162_/CLK _14162_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11374_ VGND VPWR VPWR VGND _11374_/X _14845_/Q _11392_/B _14813_/Q sky130_fd_sc_hd__mux2_1
XFILLER_4_954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10325_ VGND VPWR VPWR VGND _10325_/X hold975/A _11261_/B hold353/A sky130_fd_sc_hd__mux2_1
XFILLER_3_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10256_ VGND VPWR VGND VPWR _10256_/X _10930_/C1 _10255_/X _10252_/X _12869_/A1 sky130_fd_sc_hd__o211a_1
X_10187_ VPWR VGND VGND VPWR _10187_/X _10705_/A _10187_/B sky130_fd_sc_hd__or2_1
XFILLER_19_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14995_ hold263/A _14995_/CLK _14995_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_58_clk clkload37/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_13042__159 VPWR VGND VPWR VGND _14285_/CLK clkload24/A sky130_fd_sc_hd__inv_2
XFILLER_35_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15616_ _15616_/Q clkload27/A _15616_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12828_ VPWR VGND VGND VPWR _12826_/Y _12827_/Y _15564_/Q _10056_/A _15564_/D _07544_/B
+ sky130_fd_sc_hd__o221a_1
X_15547_ _15547_/Q clkload43/A _15547_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12759_ VPWR VGND VGND VPWR _12829_/S _08218_/Y _08222_/X _12789_/A _12759_/X _12807_/A1
+ sky130_fd_sc_hd__o221a_1
XFILLER_43_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15478_ _15478_/Q _15478_/CLK _15478_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_574 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14429_ hold947/A _14429_/CLK _14429_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold715 hold715/X hold715/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout8 VPWR VGND fanout8/X fanout9/A VPWR VGND sky130_fd_sc_hd__buf_2
Xhold726 hold726/X hold726/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 hold737/X hold737/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold704 hold704/X hold704/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ VPWR VGND VGND VPWR _09970_/A _09970_/B _09970_/Y sky130_fd_sc_hd__nor2_1
X_13740__857 VPWR VGND VPWR VGND _15112_/CLK clkload46/A sky130_fd_sc_hd__inv_2
Xhold748 hold748/X hold748/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 hold759/X hold759/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08921_ VGND VPWR VGND VPWR _15132_/D hold1115/X _08902_/B _08920_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
X_08852_ VGND VPWR _15262_/Q _08853_/B _15263_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07803_ VPWR VGND VGND VPWR _07803_/A _07909_/B _07803_/B sky130_fd_sc_hd__nand2_1
Xhold1404 hold1404/X _14843_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 hold1415/X _15066_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 hold1437/X _15696_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _08476_/A _15338_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13593__710 VPWR VGND VPWR VGND _14924_/CLK clkload54/A sky130_fd_sc_hd__inv_2
Xhold1426 hold1426/X _15089_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1448 hold1448/X _15297_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_49_clk clkload41/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_08783_ _15226_/D fanout92/X fanout88/X _08781_/Y _08782_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07734_ VPWR VGND VGND VPWR _07795_/C _15557_/Q _07734_/B sky130_fd_sc_hd__or2_1
XFILLER_38_663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_53_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07665_ VPWR VGND VGND VPWR _07665_/C _07665_/B _07665_/A _07665_/Y sky130_fd_sc_hd__nor3_1
X_09404_ VGND VPWR VPWR VGND _14645_/D hold607/X _09414_/S fanout8/X sky130_fd_sc_hd__mux2_1
X_13634__751 VPWR VGND VPWR VGND _14974_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_07596_ VGND VPWR VGND VPWR _07570_/X _08214_/A _08151_/B _07595_/Y _07596_/X sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09335_ VGND VPWR VPWR VGND _14709_/D hold572/X _09345_/S fanout10/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09266_ VGND VPWR VPWR VGND _14777_/D fanout7/X _09268_/S hold357/X sky130_fd_sc_hd__mux2_1
X_08217_ VPWR VGND VGND VPWR _08173_/Y _08216_/X _08172_/X _10583_/A2 _08217_/X _10058_/A1
+ sky130_fd_sc_hd__o221a_1
X_09197_ VGND VPWR VPWR VGND _14894_/D hold369/X _09197_/S fanout97/X sky130_fd_sc_hd__mux2_1
X_08148_ VPWR VGND VPWR VGND _15614_/Q _08299_/A2 _08148_/X _12833_/A _08145_/Y _08147_/Y
+ sky130_fd_sc_hd__a221o_1
X_08079_ VPWR VGND VPWR VGND _08100_/B _08102_/A _07195_/A _08080_/B sky130_fd_sc_hd__a21oi_1
X_11090_ VGND VPWR VPWR VGND _11090_/X _14214_/Q _11093_/S _15222_/Q sky130_fd_sc_hd__mux2_1
X_10110_ VPWR VGND VGND VPWR _10110_/X hold214/A _10521_/B sky130_fd_sc_hd__or2_1
X_10041_ VPWR VGND _10045_/C _10042_/B _15633_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_27_1424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13889__1006 VPWR VGND VPWR VGND _15261_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_14780_ hold854/A _14780_/CLK _14780_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11992_ VPWR VGND VGND VPWR _12103_/A _11992_/B _11992_/Y sky130_fd_sc_hd__nor2_1
X_10943_ VGND VPWR VPWR VGND _10943_/X hold552/A _11167_/S hold339/A sky130_fd_sc_hd__mux2_1
XFILLER_45_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13377__494 VPWR VGND VPWR VGND _14652_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_10874_ VGND VPWR VGND VPWR _10874_/X _10871_/X _10873_/X _10890_/A _10891_/C1 sky130_fd_sc_hd__a211o_1
Xclkbuf_3_0_0_clk clkbuf_3_0_0_clk/X clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12613_ VGND VPWR VPWR VGND _12613_/X _14279_/Q _12635_/B _14311_/Q sky130_fd_sc_hd__mux2_1
X_15401_ hold530/A _15401_/CLK _15401_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15332_ _15332_/Q _15332_/CLK _15332_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_40_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12544_ VGND VPWR VPWR VGND _12544_/X _12541_/X _12665_/S _12540_/X sky130_fd_sc_hd__mux2_1
X_14060__1177 VPWR VGND VPWR VGND _15479_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_15263_ _15263_/Q _15263_/CLK _15263_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_8_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12475_ VGND VPWR VPWR VGND _12475_/X hold776/A _12479_/S hold446/A sky130_fd_sc_hd__mux2_1
X_11426_ VGND VPWR VGND VPWR _11426_/X _14928_/Q _11303_/A _11431_/A2 sky130_fd_sc_hd__a21bo_1
X_14214_ _14214_/Q _14214_/CLK _14214_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_6 _07690_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_15194_ _15194_/Q _15194_/CLK _15194_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14145_ hold149/A _14145_/CLK _14145_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11357_ VPWR VGND VGND VPWR _11408_/B _14856_/Q _14855_/Q sky130_fd_sc_hd__or2_1
X_10308_ VPWR VGND VGND VPWR _10308_/X hold279/A _11098_/S sky130_fd_sc_hd__or2_1
X_11288_ VPWR VGND _14812_/D _11288_/B _11290_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_10239_ VGND VPWR VPWR VGND _10243_/B hold753/A _10258_/B hold347/A sky130_fd_sc_hd__mux2_1
XFILLER_55_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13618__735 VPWR VGND VPWR VGND _14958_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
Xrebuffer29 VPWR VGND VPWR VGND rebuffer29/X rebuffer30/X sky130_fd_sc_hd__dlygate4sd1_1
X_14978_ hold343/A _14978_/CLK _14978_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07450_ VPWR VGND VGND VPWR _07452_/B _07450_/A _07450_/B sky130_fd_sc_hd__or2_1
X_07381_ VGND VPWR VGND VPWR _07380_/X _07088_/Y _07258_/B _07381_/X sky130_fd_sc_hd__o21ba_1
X_09120_ VGND VPWR VPWR VGND _14975_/D hold412/X _09128_/S _09547_/A1 sky130_fd_sc_hd__mux2_1
XFILLER_31_850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09051_ VGND VPWR VPWR VGND _15039_/D hold616/X _09051_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
X_13170__287 VPWR VGND VPWR VGND _14445_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_08002_ VPWR VGND VPWR VGND _15621_/Q _08002_/A2 _08014_/B _08002_/B1 _15585_/Q _08001_/Y
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold501 hold501/X hold501/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 hold545/X hold545/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 hold512/X hold512/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/X hold534/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 hold523/X hold523/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 hold567/X hold567/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 hold578/X hold578/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 hold556/X hold556/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ VGND VPWR _09954_/C _09954_/B _09953_/Y _14127_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold589 hold589/X hold589/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09884_ VPWR VGND VGND VPWR hold1172/X _09880_/Y _09883_/Y _09884_/X sky130_fd_sc_hd__o21a_1
X_08904_ VPWR VGND VGND VPWR _08904_/X _15140_/Q _08924_/B sky130_fd_sc_hd__or2_1
Xhold1212 hold1212/X _14889_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 hold1234/X _14622_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1223 hold1223/X _14796_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ VGND VPWR VPWR VGND _15178_/D _08014_/X _08842_/S hold393/X sky130_fd_sc_hd__mux2_1
Xhold1201 hold1201/X _14745_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _14841_/D _11354_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 hold1245/X _15393_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 hold1267/X _15508_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ VGND VPWR VPWR VGND _15240_/D fanout20/X _08776_/S hold220/X sky130_fd_sc_hd__mux2_1
X_13064__181 VPWR VGND VPWR VGND _14307_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_07717_ VPWR VGND VGND VPWR _15562_/Q _07717_/B _07718_/B sky130_fd_sc_hd__nor2_1
Xhold1278 hold1278/X _15623_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 _10014_/A _15621_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08697_ VGND VPWR VGND VPWR _08697_/X _08700_/A2 _08700_/B1 hold1441/X _08696_/X
+ sky130_fd_sc_hd__a211o_1
X_07648_ VPWR VGND VPWR VGND _07663_/B _07663_/A _07665_/A _07664_/A sky130_fd_sc_hd__a21oi_1
X_07579_ VGND VPWR VPWR VGND _09010_/B _15546_/Q _08591_/B _10060_/C _07578_/Y sky130_fd_sc_hd__o2bb2a_1
X_09318_ VGND VPWR VPWR VGND _14726_/D _09342_/S hold1132/X clone111/X sky130_fd_sc_hd__mux2_4
X_13411__528 VPWR VGND VPWR VGND _14686_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_16_1158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10590_ VGND VPWR VPWR VGND _10590_/X hold712/A _10742_/S hold238/A sky130_fd_sc_hd__mux2_1
X_09249_ VGND VPWR VPWR VGND _14794_/D fanout70/X _09269_/S hold641/X sky130_fd_sc_hd__mux2_1
X_12260_ VGND VPWR VPWR VGND _12260_/X hold599/A _12339_/B hold206/A sky130_fd_sc_hd__mux2_1
X_12191_ VPWR VGND VGND VPWR _12191_/X hold419/A _12191_/B sky130_fd_sc_hd__or2_1
X_11211_ VGND VPWR VPWR VGND _11211_/X hold934/A _11216_/S hold709/A sky130_fd_sc_hd__mux2_1
X_11142_ VGND VPWR VPWR VGND _11142_/X hold793/A _11142_/S hold598/A sky130_fd_sc_hd__mux2_1
X_11073_ VGND VPWR VGND VPWR _11073_/X _15507_/Q _11252_/A2 _11072_/X _11250_/S sky130_fd_sc_hd__o211a_1
X_13305__422 VPWR VGND VPWR VGND _14580_/CLK clkload18/A sky130_fd_sc_hd__inv_2
XFILLER_76_522 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10024_ VGND VPWR _10028_/B _15626_/Q _15625_/Q _10024_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14901_ hold411/A _14901_/CLK _14901_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14832_ _14832_/Q _14832_/CLK _14832_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_599 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_57_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_40_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14763_ _14763_/Q _14763_/CLK _14763_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11975_ VGND VPWR VPWR VGND _11979_/B hold916/A _12005_/S hold632/A sky130_fd_sc_hd__mux2_1
X_14694_ hold570/A _14694_/CLK _14694_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_912 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10926_ VGND VPWR VGND VPWR _10926_/X _10923_/X _10925_/X _11189_/A1 _11254_/C1 sky130_fd_sc_hd__a211o_1
X_10857_ VPWR VGND VPWR VGND _10857_/X _11173_/A _10830_/X _10838_/X _10856_/X _10855_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_32_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_73_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10788_ VGND VPWR VPWR VGND _10788_/X _10787_/X _11213_/S _10786_/X sky130_fd_sc_hd__mux2_1
X_15315_ _15315_/Q _15315_/CLK _15315_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12527_ VPWR VGND _12527_/X _12526_/X _12522_/X _12731_/S _12518_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15246_ hold321/A _15246_/CLK _15246_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12458_ VGND VPWR VPWR VGND _12458_/X hold482/A _12479_/S hold313/A sky130_fd_sc_hd__mux2_1
X_11409_ VPWR VGND VGND VPWR _11406_/X _11408_/X _08541_/A _14856_/D sky130_fd_sc_hd__o21a_1
X_15177_ hold407/A _15177_/CLK _15177_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12389_ VPWR VGND VPWR VGND _12388_/X _12415_/C1 _12387_/X _12389_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14128_ _14128_/Q _14128_/CLK _14128_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Right_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13048__165 VPWR VGND VPWR VGND _14291_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
XFILLER_80_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08620_ VPWR VGND VGND VPWR _08626_/A _09013_/B _08620_/Y sky130_fd_sc_hd__nor2_1
X_13852__969 VPWR VGND VPWR VGND _15224_/CLK clkload41/A sky130_fd_sc_hd__inv_2
XFILLER_78_1141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08551_ VPWR VGND VGND VPWR _08605_/A _08974_/B _08551_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08482_ VPWR VGND VGND VPWR _08482_/X _15335_/Q _08482_/B sky130_fd_sc_hd__or2_1
X_07502_ VPWR VGND VGND VPWR _07503_/B _15463_/Q _07507_/B sky130_fd_sc_hd__or2_1
X_07433_ VPWR VGND VGND VPWR _07433_/A _07433_/B _07551_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_956 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_39_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Right_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07364_ VPWR VGND VPWR VGND _07366_/A _07222_/B _07222_/A _10062_/A _07234_/A _07234_/B
+ sky130_fd_sc_hd__o32a_1
X_09103_ VGND VPWR VPWR VGND _14992_/D hold358/X _09124_/S fanout64/X sky130_fd_sc_hd__mux2_1
X_13746__863 VPWR VGND VPWR VGND _15118_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_07295_ VPWR VGND _07298_/A _07297_/B _15467_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_13888__1005 VPWR VGND VPWR VGND _15260_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_09034_ VGND VPWR VPWR VGND _15056_/D hold527/X _09055_/S fanout64/X sky130_fd_sc_hd__mux2_1
Xhold320 hold320/X hold320/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/X hold353/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 hold342/X hold342/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 hold331/X hold331/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_518 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_77_17 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout800 VPWR VGND _08605_/A _08562_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xhold364 hold364/X hold364/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 hold386/X hold386/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold375/X hold375/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout833 VPWR VGND _09000_/C1 _09017_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout811 VPWR VGND _08735_/C fanout829/X VPWR VGND sky130_fd_sc_hd__buf_4
X_09936_ VPWR VGND _14763_/D _08425_/A _15365_/Q _14767_/Q _09938_/A VGND VPWR sky130_fd_sc_hd__a31o_1
Xfanout822 VPWR VGND _11315_/A1 fanout824/X VPWR VGND sky130_fd_sc_hd__buf_2
Xhold397 hold397/X hold397/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout844 VGND VPWR _14154_/Q fanout844/X VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout866 VPWR VGND _11303_/A _07109_/Y VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_58_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout855 VPWR VGND _07857_/A _07984_/S VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_24_1405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1031 hold1031/X _15106_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout877 VPWR VGND _09311_/B _15580_/Q VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout888 VPWR VGND _10056_/A _14802_/Q VPWR VGND sky130_fd_sc_hd__buf_4
Xhold1020 hold1020/X _15269_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 hold1042/X _14363_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09867_ VGND VPWR VPWR VGND _14155_/D hold625/X _09867_/S fanout95/X sky130_fd_sc_hd__mux2_1
Xhold1075 hold1075/X _15315_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1053 hold1053/X _15020_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ VPWR VGND VGND VPWR _08818_/X _08818_/A _08846_/S sky130_fd_sc_hd__or2_1
X_09798_ VGND VPWR VPWR VGND _14251_/D fanout97/X _09798_/S hold366/X sky130_fd_sc_hd__mux2_1
Xhold1064 hold1064/X _15504_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 hold1097/X _15103_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ VGND VPWR VPWR VGND _15257_/D fanout84/X _08773_/S hold553/X sky130_fd_sc_hd__mux2_1
XFILLER_2_1234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1086 hold1086/X _14999_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_1214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11760_ VPWR VGND VPWR VGND _11759_/X _12101_/A1 _11758_/X _11760_/Y sky130_fd_sc_hd__a21oi_1
X_10711_ VGND VPWR VGND VPWR _14395_/D _12121_/B1 _10709_/X _10710_/X _11290_/A sky130_fd_sc_hd__o211a_1
X_11691_ VPWR VGND VGND VPWR _11691_/X _12476_/S _11691_/B sky130_fd_sc_hd__or2_1
XFILLER_70_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10642_ VPWR VGND VGND VPWR _10642_/X _10652_/S _10642_/B sky130_fd_sc_hd__or2_1
X_10573_ VGND VPWR VPWR VGND _10573_/X hold383/A _10730_/S hold514/A sky130_fd_sc_hd__mux2_1
X_15100_ _15100_/Q _15100_/CLK _15100_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12312_ VPWR VGND VGND VPWR _12312_/X _12581_/S _12312_/B sky130_fd_sc_hd__or2_1
Xrebuffer9 VPWR VGND VPWR VGND _07143_/A1 _07826_/A sky130_fd_sc_hd__dlygate4sd1_1
X_12243_ VGND VPWR VPWR VGND _12243_/X hold867/A _12318_/S hold508/A sky130_fd_sc_hd__mux2_1
X_15031_ hold892/A _15031_/CLK _15031_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_378 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12174_ VGND VPWR VPWR VGND _12174_/X _12171_/X _12174_/S _12170_/X sky130_fd_sc_hd__mux2_1
X_11125_ VGND VPWR VPWR VGND _11125_/X _11122_/X _11143_/S _11121_/X sky130_fd_sc_hd__mux2_1
X_11056_ VGND VPWR VPWR VGND _11056_/X hold658/A _11165_/S hold296/A sky130_fd_sc_hd__mux2_1
XFILLER_1_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10007_ VPWR VGND VGND VPWR _10007_/A _10007_/B _10008_/B sky130_fd_sc_hd__nor2_1
XFILLER_77_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14815_ _14815_/Q clkload20/A _14815_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13689__806 VPWR VGND VPWR VGND _15029_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_14746_ hold193/A _14746_/CLK _14746_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11958_ VPWR VGND VGND VPWR _11958_/X _11958_/A _11958_/B sky130_fd_sc_hd__or2_1
XFILLER_75_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14677_ hold849/A _14677_/CLK _14677_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11889_ VGND VPWR VPWR VGND _11889_/X _15007_/Q _12191_/B hold412/A sky130_fd_sc_hd__mux2_1
X_10909_ VPWR VGND VGND VPWR _10909_/X _10911_/S _10909_/B sky130_fd_sc_hd__or2_1
X_13433__550 VPWR VGND VPWR VGND _14708_/CLK clkload17/A sky130_fd_sc_hd__inv_2
XFILLER_13_680 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15229_ hold215/A _15229_/CLK _15229_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout107 VGND VPWR _12829_/S _12820_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_47_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout129 VGND VPWR _09548_/A1 _09860_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07982_ VPWR VGND VGND VPWR _07983_/B _07982_/B _08007_/A _07981_/A sky130_fd_sc_hd__nand3b_1
Xfanout118 VGND VPWR _09655_/A0 _09829_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_13282__399 VPWR VGND VPWR VGND _14557_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_09721_ VGND VPWR VPWR VGND _14322_/D _09860_/A0 _09721_/S hold761/X sky130_fd_sc_hd__mux2_1
X_09652_ VGND VPWR VPWR VGND _14418_/D hold919/X _09659_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_08603_ VGND VPWR _08603_/B _08603_/Y _08603_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_09583_ VGND VPWR VPWR VGND _14482_/D hold969/X _09590_/S _09860_/A0 sky130_fd_sc_hd__mux2_1
X_08534_ VPWR VGND VPWR VGND _08534_/B1 _15318_/Q _08540_/A2 _08535_/B _15319_/Q sky130_fd_sc_hd__a22o_1
Xtt_um_femto_889 uio_oe[0] tt_um_femto_889/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_63_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08465_ VGND VPWR VGND VPWR _08465_/X hold1290/X _08483_/A2 _08464_/X _11974_/C1
+ sky130_fd_sc_hd__o211a_1
X_13176__293 VPWR VGND VPWR VGND _14451_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_07416_ VPWR VGND VGND VPWR _07416_/A _10075_/A _07416_/Y sky130_fd_sc_hd__nor2_1
X_08396_ VGND VPWR VPWR VGND _15381_/D fanout28/X _08411_/S hold756/X sky130_fd_sc_hd__mux2_1
X_07347_ _07347_/X _07280_/B _15464_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_09017_ VPWR VGND _15098_/D _09017_/B _09017_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07278_ VPWR VGND VGND VPWR _15464_/Q _07280_/B _07926_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold150 hold150/X hold150/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 hold161/X hold161/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/X hold183/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold172/X hold172/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/X hold194/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 _09760_/S _09729_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_59_820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout641 VPWR VGND _09588_/S _09557_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_09919_ VPWR VGND VGND VPWR _14140_/Q _09923_/D _09931_/B _09919_/Y sky130_fd_sc_hd__nor3_2
Xfanout652 _09517_/S _09486_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout663 _09304_/S _09307_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout685 VPWR VGND _08356_/S _08372_/S VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_8_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout674 VGND VPWR _09095_/X _09126_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout696 VGND VPWR _08926_/B _08924_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_13874__991 VPWR VGND VPWR VGND _15246_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_73_322 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12861_ VGND VPWR VPWR VGND _15585_/D _12861_/A1 _12870_/S hold1325/X sky130_fd_sc_hd__mux2_1
X_11812_ VGND VPWR VGND VPWR _11812_/X hold975/A _12746_/A2 _12748_/A1 _11811_/X sky130_fd_sc_hd__o211a_1
XFILLER_46_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14600_ hold403/A _14600_/CLK _14600_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15580_ _15580_/Q clkload31/A _15580_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12792_ VPWR VGND VGND VPWR _10078_/A _12833_/B _08037_/Y _12792_/X sky130_fd_sc_hd__o21a_1
X_13417__534 VPWR VGND VPWR VGND _14692_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_11743_ VPWR VGND VGND VPWR _11743_/X hold327/A _12726_/S sky130_fd_sc_hd__or2_1
X_14531_ hold179/A _14531_/CLK _14531_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11674_ VGND VPWR VGND VPWR _11674_/X _15001_/Q _12192_/A2 _12180_/S _11673_/X sky130_fd_sc_hd__o211a_1
X_14462_ hold378/A _14462_/CLK _14462_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10625_ VGND VPWR VPWR VGND _10625_/X _10624_/X _10625_/S _10623_/X sky130_fd_sc_hd__mux2_1
X_14393_ _14393_/Q clkload7/A _14393_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_6_610 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10556_ VGND VPWR VGND VPWR _10556_/X _10557_/A _10552_/X _10555_/X _10717_/C1 sky130_fd_sc_hd__o211a_1
X_10487_ VPWR VGND _10487_/X _10486_/X _10482_/X _10469_/S _10478_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12975__92 VPWR VGND VPWR VGND _14218_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_13959__1076 VPWR VGND VPWR VGND _15331_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_15014_ _15014_/Q _15014_/CLK _15014_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12226_ VGND VPWR VGND VPWR _12226_/X _12223_/X _12225_/X _12226_/A1 _12226_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_69_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12984__101 VPWR VGND VPWR VGND _14227_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_12157_ VPWR VGND _12157_/X _12156_/X _12152_/X _12139_/S _12148_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11108_ VGND VPWR VPWR VGND _11112_/B _15508_/Q _11109_/S _14534_/Q sky130_fd_sc_hd__mux2_1
X_12088_ VGND VPWR VPWR VGND _12088_/X hold451/A _12097_/S hold593/A sky130_fd_sc_hd__mux2_1
XFILLER_49_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11039_ VGND VPWR VGND VPWR _11039_/X hold914/A _11184_/A2 _11038_/X _11250_/S sky130_fd_sc_hd__o211a_1
X_13887__1004 VPWR VGND VPWR VGND _15259_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14729_ hold911/A _14729_/CLK _14729_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08250_ VGND VPWR VGND VPWR _08248_/X _08250_/X _08250_/A _08250_/B sky130_fd_sc_hd__or3b_4
X_08181_ VPWR VGND _08181_/X _08181_/B _08181_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07201_ VPWR VGND _08115_/A _07358_/B _15453_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07132_ VPWR VGND VGND VPWR _09799_/A _08377_/A _07132_/Y sky130_fd_sc_hd__nor2_1
X_13210__327 VPWR VGND VPWR VGND _14485_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_13858__975 VPWR VGND VPWR VGND _15230_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_07965_ VGND VPWR _07965_/B _12810_/B _07971_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_68_683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09704_ VGND VPWR VPWR VGND _14339_/D fanout61/X _09725_/S hold482/X sky130_fd_sc_hd__mux2_1
X_07896_ VGND VPWR _07811_/B _07899_/A _07897_/B _07811_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_13104__221 VPWR VGND VPWR VGND _14347_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_09635_ VGND VPWR VPWR VGND _14435_/D hold939/X _09656_/S fanout62/X sky130_fd_sc_hd__mux2_1
XFILLER_36_580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09566_ VGND VPWR VPWR VGND _14499_/D hold1039/X _09587_/S fanout61/X sky130_fd_sc_hd__mux2_1
X_08517_ VPWR VGND VPWR VGND _08534_/B1 hold1416/X _08503_/A _08518_/B hold1418/X
+ sky130_fd_sc_hd__a22o_1
X_09497_ VGND VPWR VPWR VGND _14562_/D fanout58/X _09514_/S hold603/X sky130_fd_sc_hd__mux2_1
X_08448_ VPWR VGND VGND VPWR _08448_/A _08448_/Y _08448_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_263 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10410_ VPWR VGND VGND VPWR _10410_/X hold412/A _10702_/S sky130_fd_sc_hd__or2_1
X_08379_ VPWR VGND VGND VPWR _08379_/X _08379_/A _08405_/S sky130_fd_sc_hd__or2_1
XFILLER_11_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11390_ VGND VPWR VGND VPWR _11390_/X _14850_/Q _11362_/X _11389_/X _11388_/S sky130_fd_sc_hd__o211a_1
XFILLER_20_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10341_ VGND VPWR VGND VPWR _14385_/D _12602_/B1 _10339_/X _10340_/X _11341_/A sky130_fd_sc_hd__o211a_1
XFILLER_3_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10272_ VPWR VGND VGND VPWR _10272_/X _10613_/A _10272_/B sky130_fd_sc_hd__or2_1
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12011_ VPWR VGND VGND VPWR _11992_/Y _12010_/X _10192_/B _15456_/Q _15456_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout493 VPWR VGND _11954_/S fanout497/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout460 VGND VPWR clone2/A _11209_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout471 VPWR VGND _12669_/A2 _12080_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout482 VGND VPWR _12006_/B _11998_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_15701_ VGND VPWR _15701_/A uo_out[6] VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15632_ _15632_/Q clkload49/A _15632_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_34_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12844_ VPWR VGND VGND VPWR _12842_/X _12843_/X _11477_/S _15570_/D sky130_fd_sc_hd__o21a_1
XFILLER_76_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12775_ VGND VPWR VPWR VGND _15551_/D _12774_/X _12773_/X _12807_/A1 _12807_/B1 _15551_/Q
+ sky130_fd_sc_hd__a32o_1
X_15563_ _15563_/Q clkload44/A _15563_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13651__768 VPWR VGND VPWR VGND _14991_/CLK clkload37/A sky130_fd_sc_hd__inv_2
XFILLER_37_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14514_ hold194/A _14514_/CLK _14514_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11726_ VGND VPWR VPWR VGND _11726_/X _14191_/Q _11748_/S hold264/A sky130_fd_sc_hd__mux2_1
XFILLER_14_285 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15494_ _15494_/Q _15494_/CLK _15494_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14445_ hold681/A _14445_/CLK _14445_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11657_ VPWR VGND VPWR VGND _11656_/X _12185_/A1 _11655_/X _11657_/Y sky130_fd_sc_hd__a21oi_1
X_11588_ VGND VPWR VPWR VGND _11588_/X _11587_/X _11625_/S _11586_/X sky130_fd_sc_hd__mux2_1
X_10608_ VPWR VGND VPWR VGND _10607_/X _10608_/A1 _10606_/X _10608_/Y sky130_fd_sc_hd__a21oi_1
X_14376_ _14376_/Q _14376_/CLK _14376_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold908 hold908/X hold908/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ VPWR VGND VGND VPWR _10539_/X hold227/A _10700_/S sky130_fd_sc_hd__or2_1
Xhold919 hold919/X hold919/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13545__662 VPWR VGND VPWR VGND _14876_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_12209_ VPWR VGND VGND VPWR _12209_/X _12221_/S _12209_/B sky130_fd_sc_hd__or2_1
XFILLER_78_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07750_ _08146_/A _07748_/X _07750_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_65_642 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07681_ VPWR VGND VGND VPWR _07681_/Y _07681_/B _07681_/C _07665_/B sky130_fd_sc_hd__nand3b_1
XFILLER_20_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09420_ VGND VPWR VPWR VGND _09443_/S fanout81/X hold1191/X _14632_/D sky130_fd_sc_hd__mux2_2
X_09351_ VGND VPWR VPWR VGND _14695_/D hold487/X _09357_/S clone146/X sky130_fd_sc_hd__mux2_1
X_08302_ VGND VPWR VGND VPWR _15580_/Q _12855_/A0 _15639_/Q _15581_/Q _09521_/A sky130_fd_sc_hd__and4bb_1
X_09282_ VGND VPWR VPWR VGND _14759_/D fanout78/X _09304_/S hold287/X sky130_fd_sc_hd__mux2_1
X_08233_ VPWR VGND VGND VPWR _08233_/X _08233_/A _08233_/B sky130_fd_sc_hd__or2_1
X_08164_ VGND VPWR VGND VPWR _08164_/X _08162_/Y _08163_/X _08280_/B2 _08157_/Y sky130_fd_sc_hd__o211a_1
X_07115_ VPWR VGND VPWR VGND _08505_/A _09912_/A sky130_fd_sc_hd__inv_2
X_08095_ VPWR VGND VGND VPWR _08094_/X _07421_/Y _08093_/X _07421_/A _08095_/X _07996_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_47_1054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14029__1146 VPWR VGND VPWR VGND _15401_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XFILLER_76_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08997_ VGND VPWR VGND VPWR _15105_/D hold904/X _09015_/A2 _08996_/X _11347_/A sky130_fd_sc_hd__o211a_1
XFILLER_5_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07948_ _07953_/B _07944_/X _07945_/Y _07947_/X _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_5_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07879_ VGND VPWR VPWR VGND _07879_/X _07878_/X _07984_/S _12826_/B sky130_fd_sc_hd__mux2_1
X_10890_ VPWR VGND VGND VPWR _10890_/X _10890_/A _10890_/B sky130_fd_sc_hd__or2_1
X_09618_ VGND VPWR VPWR VGND _14450_/D _09826_/A1 _09625_/S hold1089/X sky130_fd_sc_hd__mux2_1
X_13958__1075 VPWR VGND VPWR VGND _15330_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_09549_ VGND VPWR VPWR VGND _14513_/D _09792_/A1 _09549_/S hold286/X sky130_fd_sc_hd__mux2_1
X_13488__605 VPWR VGND VPWR VGND _14763_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_12560_ VPWR VGND VGND VPWR _12560_/X hold157/A _12671_/S sky130_fd_sc_hd__or2_1
XFILLER_11_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11511_ VGND VPWR VPWR VGND _11511_/X _15089_/Q _11535_/C _15087_/Q sky130_fd_sc_hd__mux2_1
X_12491_ VPWR VGND VPWR VGND _12490_/X _12473_/A _12491_/B1 _12491_/X sky130_fd_sc_hd__a21o_1
X_11442_ VPWR VGND VPWR VGND _11475_/S _15066_/Q _12845_/B _11442_/Y sky130_fd_sc_hd__a21oi_1
X_14230_ hold360/A _14230_/CLK _14230_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13529__646 VPWR VGND VPWR VGND _14809_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_14161_ hold551/A _14161_/CLK _14161_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11373_ VGND VPWR VPWR VGND _14844_/D _11372_/X _11382_/S hold1312/X sky130_fd_sc_hd__mux2_1
X_13886__1003 VPWR VGND VPWR VGND _15258_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_10324_ VPWR VGND VPWR VGND _10321_/X _10816_/A _10323_/X _10324_/X sky130_fd_sc_hd__a21o_1
X_12945__62 VPWR VGND VPWR VGND _14188_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_3_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_966 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10255_ VGND VPWR VPWR VGND _10255_/X _10254_/X _10911_/S _10253_/X sky130_fd_sc_hd__mux2_1
X_10186_ VGND VPWR VGND VPWR _10186_/X _10705_/A _10182_/X _10185_/X _10704_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_43_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14994_ _14994_/Q _14994_/CLK _14994_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout290 VGND VPWR _10521_/B _10516_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_35_815 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13081__198 VPWR VGND VPWR VGND _14324_/CLK clkload18/A sky130_fd_sc_hd__inv_2
XFILLER_74_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12827_ VGND VPWR _12825_/X _10056_/A _12827_/Y _12817_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_15615_ _15615_/Q clkload27/A _15615_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_50_818 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15546_ _15546_/Q clkload43/A _15546_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12758_ VPWR VGND VPWR VGND _08220_/B _10079_/X _12758_/Y _08220_/C sky130_fd_sc_hd__o21bai_1
X_15477_ _15477_/Q _15477_/CLK _15477_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12689_ VGND VPWR VPWR VGND _12689_/X hold604/A _12689_/S hold249/A sky130_fd_sc_hd__mux2_1
X_11709_ VGND VPWR VPWR VGND _11709_/X hold842/A _12716_/S hold614/A sky130_fd_sc_hd__mux2_1
X_14428_ hold798/A _14428_/CLK _14428_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout9 VPWR VGND VPWR VGND fanout9/X fanout9/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold705 hold705/X hold705/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ _14359_/Q _14359_/CLK _14359_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold727 hold727/X hold727/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 hold716/X hold716/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 hold738/X hold738/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 hold749/X hold749/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08920_ VPWR VGND VGND VPWR _08920_/X _08920_/A _08924_/B sky130_fd_sc_hd__or2_1
X_08851_ VPWR VGND VGND VPWR _09938_/A _08851_/B _15162_/D sky130_fd_sc_hd__nor2_1
XFILLER_48_1396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1416 hold1416/X _15326_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07802_ VPWR VGND VPWR VGND _07915_/B _07915_/A _07718_/A _07909_/A sky130_fd_sc_hd__a21oi_1
X_13322__439 VPWR VGND VPWR VGND _14597_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
Xhold1405 hold1405/X _15082_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1449 _09942_/A _14131_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 hold1427/X _15086_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 hold1438/X _15279_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08782_ VPWR VGND VGND VPWR _08782_/X _08782_/A _08811_/S sky130_fd_sc_hd__or2_1
X_07733_ VPWR VGND VPWR VGND _07733_/Y _07998_/B sky130_fd_sc_hd__inv_2
XFILLER_37_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_53_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07664_ VPWR VGND VGND VPWR _07664_/X _07664_/A _07664_/B sky130_fd_sc_hd__or2_1
XFILLER_38_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13673__790 VPWR VGND VPWR VGND _15013_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_09403_ VGND VPWR VPWR VGND _14646_/D hold632/X _09414_/S fanout12/X sky130_fd_sc_hd__mux2_1
X_07595_ VPWR VGND VGND VPWR _08198_/S _08232_/B _07595_/Y sky130_fd_sc_hd__nor2_1
X_09334_ VGND VPWR VPWR VGND _14710_/D hold870/X _09345_/S fanout13/X sky130_fd_sc_hd__mux2_1
X_09265_ VGND VPWR VPWR VGND _14778_/D fanout8/X _09275_/S hold879/X sky130_fd_sc_hd__mux2_1
X_13216__333 VPWR VGND VPWR VGND _14491_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_08216_ VPWR VGND VPWR VGND _08252_/A2 _15157_/Q _08215_/X _08216_/X sky130_fd_sc_hd__a21o_1
X_09196_ VGND VPWR VPWR VGND _14895_/D hold483/X _09197_/S fanout99/X sky130_fd_sc_hd__mux2_1
X_08147_ VPWR VGND VGND VPWR _08147_/A _12772_/A _08147_/Y sky130_fd_sc_hd__nor2_1
X_08078_ VPWR VGND VGND VPWR _08059_/B _08078_/B _08078_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_66_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10040_ VPWR VGND VGND VPWR _10042_/B _10040_/B _15632_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_1436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_973 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11991_ VGND VPWR VPWR VGND _11992_/B _11990_/Y _12176_/S _11982_/Y sky130_fd_sc_hd__mux2_1
XFILLER_72_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10942_ VGND VPWR VPWR VGND _10946_/B hold670/A _11167_/S hold198/A sky130_fd_sc_hd__mux2_1
XFILLER_44_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15400_ hold445/A _15400_/CLK _15400_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10873_ VGND VPWR VGND VPWR _10873_/X hold999/A _12866_/A1 _10872_/X _11110_/A sky130_fd_sc_hd__o211a_1
XFILLER_32_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12612_ VGND VPWR VPWR VGND _12616_/B _14796_/Q _12635_/B _14247_/Q sky130_fd_sc_hd__mux2_1
X_15331_ _15696_/A _15331_/CLK _15331_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12543_ VGND VPWR VGND VPWR _12543_/X _12662_/A1 _12539_/X _12542_/X _12662_/C1 sky130_fd_sc_hd__o211a_1
X_15262_ _15262_/Q _15262_/CLK _15262_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14213_ _14213_/Q _14213_/CLK _14213_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12474_ VGND VPWR VPWR VGND _12474_/X hold939/A _12479_/S hold754/A sky130_fd_sc_hd__mux2_1
X_11425_ VGND VPWR VGND VPWR _14927_/D _14928_/Q _11431_/A2 _11424_/X _11431_/C1 sky130_fd_sc_hd__o211a_1
XANTENNA_7 _07690_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_15193_ hold841/A _15193_/CLK _15193_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14144_ _14144_/Q _14144_/CLK _14144_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11356_ VPWR VGND VPWR VGND _14851_/Q _14853_/Q _14854_/Q _14852_/Q _11356_/X sky130_fd_sc_hd__or4_1
X_10307_ VGND VPWR VPWR VGND _10307_/X _10306_/X _10315_/S _10305_/X sky130_fd_sc_hd__mux2_1
X_11287_ VGND VPWR VPWR VGND _11288_/B _14812_/Q _11299_/S _14380_/Q sky130_fd_sc_hd__mux2_1
XFILLER_79_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10238_ VPWR VGND VPWR VGND _10237_/X _10930_/C1 _10236_/X _10238_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_1007 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10169_ VPWR VGND VGND VPWR _10169_/X hold278/A _10169_/B sky130_fd_sc_hd__or2_1
XFILLER_43_1260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14977_ hold391/A _14977_/CLK _14977_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13657__774 VPWR VGND VPWR VGND _14997_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_50_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07380_ _07380_/X _07252_/B _15457_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_14028__1145 VPWR VGND VPWR VGND _15400_/CLK clkload23/A sky130_fd_sc_hd__inv_2
X_15529_ hold270/A _15529_/CLK _15529_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09050_ VGND VPWR VPWR VGND _15040_/D hold696/X _09059_/S fanout5/X sky130_fd_sc_hd__mux2_1
X_08001_ VPWR VGND VGND VPWR _08147_/A _07999_/X _08000_/Y _08220_/A _08001_/Y sky130_fd_sc_hd__o22ai_1
Xhold502 hold502/X hold502/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 hold524/X hold524/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 hold513/X hold513/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 hold535/X hold535/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ VPWR VGND VPWR VGND _09951_/Y hold1383/X _09956_/S _14127_/D _09937_/Y sky130_fd_sc_hd__a22o_1
Xhold568 hold568/X hold568/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 hold557/X hold557/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 hold546/X hold546/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 hold579/X hold579/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13957__1074 VPWR VGND VPWR VGND _15329_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08903_ VGND VPWR VGND VPWR _15141_/D hold1313/X _08880_/B _08902_/Y _11399_/A1 sky130_fd_sc_hd__o211a_1
X_09883_ VPWR VGND VPWR VGND _09880_/Y _14148_/Q _09882_/A _09883_/Y sky130_fd_sc_hd__a21oi_1
Xhold1224 hold1224/X _14836_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1202 hold1202/X _14624_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ VGND VPWR VPWR VGND _15179_/D fanout33/X _08850_/S hold705/X sky130_fd_sc_hd__mux2_1
Xhold1213 hold1213/X _15280_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _08733_/A _15263_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 hold1257/X _15159_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 hold1235/X _14430_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ VGND VPWR VPWR VGND _15241_/D fanout24/X _08779_/S hold593/X sky130_fd_sc_hd__mux2_1
XFILLER_22_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_66_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1268 hold1268/X _15026_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 hold1279/X _15136_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07716_ VPWR VGND _07718_/A _07717_/B _15562_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_22_1366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13885__1002 VPWR VGND VPWR VGND _15257_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_08696_ VGND VPWR VGND VPWR _08696_/X _14393_/Q _08640_/B _08711_/B1 _08634_/X sky130_fd_sc_hd__o211a_1
XFILLER_22_1388 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07647_ VPWR VGND VPWR VGND _07908_/B1 _15633_/Q _07952_/A2 _07659_/A _15597_/Q sky130_fd_sc_hd__a22o_1
X_07578_ VGND VPWR _07578_/B _07578_/Y _07578_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13450__567 VPWR VGND VPWR VGND _14725_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_09317_ VGND VPWR VPWR VGND _14727_/D hold598/X _09327_/S fanout78/X sky130_fd_sc_hd__mux2_1
XFILLER_22_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_1137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09248_ VGND VPWR VPWR VGND _14795_/D _09269_/S clone47/A hold1231/X sky130_fd_sc_hd__mux2_4
X_09179_ VGND VPWR VPWR VGND _14912_/D hold581/X _09194_/S fanout38/X sky130_fd_sc_hd__mux2_1
X_11210_ VPWR VGND VGND VPWR _11210_/A _11210_/B _11210_/Y sky130_fd_sc_hd__nor2_1
X_12190_ VGND VPWR VPWR VGND _12190_/X hold705/A _12190_/S hold420/A sky130_fd_sc_hd__mux2_1
X_11141_ VGND VPWR VPWR VGND _11141_/X hold941/A _11146_/B hold487/A sky130_fd_sc_hd__mux2_1
X_12915__32 VPWR VGND VPWR VGND _14158_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XFILLER_27_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13344__461 VPWR VGND VPWR VGND _14619_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_11072_ VPWR VGND VGND VPWR _11072_/X hold157/A _11186_/S sky130_fd_sc_hd__or2_1
XFILLER_27_1244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14900_ hold353/A _14900_/CLK _14900_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10023_ VGND VPWR VPWR VGND _10023_/A _15625_/D _10024_/C sky130_fd_sc_hd__xor2_1
XFILLER_23_1108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14831_ _14831_/Q _14832_/CLK _14831_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_57_770 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11974_ VGND VPWR VGND VPWR _15455_/D _11974_/A1 _11972_/X _11973_/Y _11974_/C1 sky130_fd_sc_hd__o211a_1
X_14762_ _14762_/Q _14762_/CLK _14762_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14693_ hold436/A _14693_/CLK _14693_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10925_ VGND VPWR VGND VPWR _10925_/X _15503_/Q _11252_/A2 _10924_/X _11244_/S sky130_fd_sc_hd__o211a_1
XFILLER_72_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10856_ VPWR VGND _10856_/X _10846_/X _10842_/X _11218_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
X_15314_ hold942/A _15314_/CLK _15314_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10787_ VGND VPWR VPWR VGND _10787_/X _14494_/Q _11216_/S _14174_/Q sky130_fd_sc_hd__mux2_1
X_12526_ VGND VPWR VGND VPWR _12526_/X _12523_/X _12525_/X _12674_/A1 _12740_/A1 sky130_fd_sc_hd__a211o_1
X_15245_ hold182/A _15245_/CLK _15245_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12457_ VGND VPWR VPWR VGND _12457_/X _14499_/Q _12479_/S hold480/A sky130_fd_sc_hd__mux2_1
X_11408_ VGND VPWR _11408_/X _11408_/B _11408_/A _11410_/B VPWR VGND sky130_fd_sc_hd__and3_1
X_15176_ hold372/A _15176_/CLK _15176_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14127_ _14127_/Q _14127_/CLK _14127_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12388_ VGND VPWR VPWR VGND _12388_/X _12385_/X _12396_/S _12384_/X sky130_fd_sc_hd__mux2_1
X_11339_ VPWR VGND VGND VPWR _11421_/C _11316_/Y _07107_/Y _11338_/Y _11340_/B sky130_fd_sc_hd__o22a_1
XFILLER_79_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_55_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08550_ VGND VPWR VPWR VGND _08974_/B _08549_/Y _08548_/X _07534_/B _08604_/B2 _08542_/Y
+ sky130_fd_sc_hd__a32o_1
XFILLER_35_431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14208__926 _14208_/D _14208__926/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08481_ VGND VPWR VGND VPWR _15336_/D hold1198/X _08483_/A2 _08480_/X _11431_/C1
+ sky130_fd_sc_hd__o211a_1
X_07501_ VPWR VGND VGND VPWR _15463_/Q _07531_/C _07507_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_1115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_78_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07432_ VPWR VGND VGND VPWR _15461_/Q _07507_/B _07433_/B sky130_fd_sc_hd__nor2_1
X_07363_ VGND VPWR VGND VPWR _07362_/Y _07222_/B _07222_/A _08241_/B sky130_fd_sc_hd__o21ba_1
X_09102_ VGND VPWR VPWR VGND _14993_/D hold332/X _09124_/S fanout68/X sky130_fd_sc_hd__mux2_1
XFILLER_17_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_17_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07294_ VPWR VGND VGND VPWR _14401_/Q _07301_/A2 _07301_/B1 _07297_/B sky130_fd_sc_hd__o21a_1
X_09033_ VGND VPWR VPWR VGND _15057_/D hold385/X _09055_/S fanout68/X sky130_fd_sc_hd__mux2_1
X_13287__404 VPWR VGND VPWR VGND _14562_/CLK clkload42/A sky130_fd_sc_hd__inv_2
Xhold310 hold310/X hold310/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/X hold321/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold332/X hold332/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Left_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold343 hold343/X hold343/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 hold387/X hold387/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 hold354/X hold354/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 hold376/X hold376/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 hold365/X hold365/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13328__445 VPWR VGND VPWR VGND _14603_/CLK clkload12/A sky130_fd_sc_hd__inv_2
Xfanout834 VPWR VGND _11337_/C1 _09017_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout823 VPWR VGND _11431_/C1 fanout824/X VPWR VGND sky130_fd_sc_hd__buf_2
X_09935_ VPWR VGND _14132_/D _09917_/A _09934_/Y hold239/X _08498_/Y _09919_/Y VPWR
+ VGND sky130_fd_sc_hd__a311oi_1
Xfanout801 VGND VPWR fanout802/X _08562_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold398 hold398/X hold398/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout812 VPWR VGND _11294_/A _12159_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout845 VGND VPWR _11406_/C _11392_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout867 VPWR VGND _07714_/A _15601_/Q VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout856 VGND VPWR _08182_/S _07984_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09866_ VGND VPWR VPWR VGND _14156_/D hold396/X _09867_/S fanout99/X sky130_fd_sc_hd__mux2_1
Xfanout878 VGND VPWR _12855_/A0 _09556_/C VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold1010 hold1010/X _14493_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1021 hold1021/X _15396_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ VPWR VGND VPWR VGND _08817_/Y _08846_/S sky130_fd_sc_hd__inv_2
Xhold1032 hold1032/X _14422_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 hold1076/X _15102_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 hold1054/X _15304_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1065 hold1065/X _14257_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 hold1043/X _15018_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09797_ VGND VPWR VPWR VGND _14252_/D fanout98/X _09798_/S hold512/X sky130_fd_sc_hd__mux2_1
Xhold1098 _15103_/D _09003_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_1246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1087 hold1087/X _15022_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _15258_/D fanout94/X fanout90/X _08746_/Y _08747_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08679_ VPWR VGND VPWR VGND hold952/A _08562_/A _08679_/X _08691_/B1 _08678_/X _08688_/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10710_ VPWR VGND VGND VPWR _10710_/X _14395_/Q _10710_/B sky130_fd_sc_hd__or2_1
X_11690_ VGND VPWR VPWR VGND _11690_/X hold937/A _12052_/S hold423/A sky130_fd_sc_hd__mux2_1
X_10641_ VGND VPWR VPWR VGND _10641_/X hold745/A _10720_/S hold218/A sky130_fd_sc_hd__mux2_1
XFILLER_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10572_ VGND VPWR VPWR VGND _10576_/B hold574/A _10730_/S hold302/A sky130_fd_sc_hd__mux2_1
XFILLER_10_843 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12311_ VGND VPWR VPWR VGND _12311_/X hold571/A _12577_/S hold526/A sky130_fd_sc_hd__mux2_1
X_12242_ VGND VPWR VPWR VGND _12242_/X _14205_/Q _12318_/S hold277/A sky130_fd_sc_hd__mux2_1
X_15030_ _15030_/Q _15030_/CLK _15030_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_68_1388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12173_ VGND VPWR VGND VPWR _12173_/X _11958_/A _12169_/X _12172_/X _12184_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11124_ VGND VPWR VGND VPWR _11124_/X _11189_/A1 _11120_/X _11123_/X _11254_/C1 sky130_fd_sc_hd__o211a_1
X_11055_ VGND VPWR VPWR VGND _11055_/X _14213_/Q _11165_/S hold285/A sky130_fd_sc_hd__mux2_1
X_14027__1144 VPWR VGND VPWR VGND _15399_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_76_320 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10006_ VPWR VGND _10010_/C _10007_/B _15618_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_37_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14814_ _14814_/Q clkload19/A _14814_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13121__238 VPWR VGND VPWR VGND _14364_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_11957_ VGND VPWR VPWR VGND _11957_/X hold781/A _11964_/S hold699/A sky130_fd_sc_hd__mux2_1
X_14745_ _14745_/Q _14745_/CLK _14745_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10908_ VGND VPWR VPWR VGND _10908_/X _14465_/Q _10919_/S _14753_/Q sky130_fd_sc_hd__mux2_1
X_13956__1073 VPWR VGND VPWR VGND _15328_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_11888_ VGND VPWR VPWR VGND _11892_/B hold399/A _12191_/B hold616/A sky130_fd_sc_hd__mux2_1
X_14676_ hold836/A _14676_/CLK _14676_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13769__886 VPWR VGND VPWR VGND _15141_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_10839_ VGND VPWR VPWR VGND _10839_/X hold785/A _10850_/S hold565/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_34_1078 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12509_ VGND VPWR VPWR VGND _12510_/B _12508_/Y _12731_/S _12500_/Y sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13015__132 VPWR VGND VPWR VGND _14258_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_15228_ hold318/A _15228_/CLK _15228_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13884__1001 VPWR VGND VPWR VGND _15256_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_15159_ _15159_/Q _15159_/CLK _15159_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout108 VGND VPWR _10078_/Y _12829_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_07981_ VGND VPWR _07981_/B _12806_/B _07981_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xfanout119 VGND VPWR _09655_/A0 _09689_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09720_ VGND VPWR VPWR VGND _14323_/D _09825_/A1 _09728_/S hold884/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09651_ VGND VPWR VPWR VGND _14419_/D hold933/X _09659_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
X_08602_ VGND VPWR VGND VPWR _15307_/D hold1122/X _08613_/A2 _08601_/X _09000_/C1
+ sky130_fd_sc_hd__o211a_1
X_09582_ VGND VPWR VPWR VGND _14483_/D hold1090/X _09590_/S _09859_/A0 sky130_fd_sc_hd__mux2_1
X_08533_ VPWR VGND _15320_/D _08533_/B _11398_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_13713__830 VPWR VGND VPWR VGND _15053_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_70_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08464_ VPWR VGND VGND VPWR _08464_/X _15344_/Q _08482_/B sky130_fd_sc_hd__or2_1
XFILLER_51_743 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_56_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07415_ VPWR VGND VGND VPWR _15584_/Q _07415_/Y _07574_/A sky130_fd_sc_hd__nand2_1
X_08395_ VGND VPWR VPWR VGND _15382_/D fanout34/X _08411_/S hold528/X sky130_fd_sc_hd__mux2_1
XFILLER_17_1210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_50_297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07346_ VPWR VGND VPWR VGND _07180_/B _15462_/Q _07345_/X _07942_/B sky130_fd_sc_hd__a21o_1
X_09016_ VPWR VGND VPWR VGND _09016_/B1 hold1443/X _08933_/A _09017_/B _15098_/Q sky130_fd_sc_hd__a22o_1
X_07277_ VPWR VGND VGND VPWR _14398_/Q _07304_/A2 _07304_/B1 _07280_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold151 hold151/X hold151/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13562__679 VPWR VGND VPWR VGND _14893_/CLK clkload39/A sky130_fd_sc_hd__inv_2
Xhold162 hold162/X hold162/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/X hold173/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/X hold195/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/X hold184/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout642 _09584_/S _09587_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09918_ VPWR VGND VGND VPWR _14138_/Q _09916_/B hold1371/X _09918_/X sky130_fd_sc_hd__o21a_1
Xfanout631 VPWR VGND _09693_/S _09684_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout620 VPWR VGND _09865_/S _09834_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout664 _09307_/S _09276_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout675 VPWR VGND _09124_/S _09125_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout653 _09485_/S _09478_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout697 VGND VPWR _08918_/B _08926_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09849_ VGND VPWR VPWR VGND _14173_/D hold855/X _09861_/S fanout40/X sky130_fd_sc_hd__mux2_1
Xfanout686 _08372_/S _08342_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12860_ VGND VPWR VPWR VGND _15584_/D _08016_/X _12860_/S _15584_/Q sky130_fd_sc_hd__mux2_1
XFILLER_61_518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11811_ VPWR VGND VGND VPWR _11811_/X hold353/A _12747_/S sky130_fd_sc_hd__or2_1
XFILLER_37_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12791_ VGND VPWR VPWR VGND _15555_/D _12790_/Y _12789_/Y _12807_/A1 _12807_/B1 _15555_/Q
+ sky130_fd_sc_hd__a32o_1
X_13456__573 VPWR VGND VPWR VGND _14731_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_14530_ hold156/A _14530_/CLK _14530_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11742_ VGND VPWR VPWR VGND _11742_/X hold609/A _12726_/S hold768/A sky130_fd_sc_hd__mux2_1
X_11673_ VPWR VGND VGND VPWR _11673_/X hold777/A _11965_/S sky130_fd_sc_hd__or2_1
X_14461_ hold867/A _14461_/CLK _14461_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_916 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10624_ VGND VPWR VPWR VGND _10624_/X hold949/A _10632_/B hold724/A sky130_fd_sc_hd__mux2_1
X_14392_ _14392_/Q clkload16/A _14392_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10555_ VPWR VGND VGND VPWR _10555_/X _10662_/S _10555_/B sky130_fd_sc_hd__or2_1
X_10486_ VGND VPWR VGND VPWR _10486_/X _10483_/X _10485_/X _10486_/A1 _10693_/B1 sky130_fd_sc_hd__a211o_1
X_15013_ _15013_/Q _15013_/CLK _15013_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12225_ VGND VPWR VGND VPWR _12225_/X hold926/A _12229_/A2 _12069_/S _12224_/X sky130_fd_sc_hd__o211a_1
X_12156_ VGND VPWR VGND VPWR _12156_/X _12155_/X _12154_/X _12156_/A1 _12202_/C1 sky130_fd_sc_hd__a211o_1
X_11107_ VGND VPWR VPWR VGND _11107_/X _15026_/Q _11107_/S _14994_/Q sky130_fd_sc_hd__mux2_1
XFILLER_1_371 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_42_1325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12087_ VGND VPWR VPWR VGND _12087_/X _14489_/Q _12094_/S hold351/A sky130_fd_sc_hd__mux2_1
X_11038_ VPWR VGND VGND VPWR _11038_/X hold295/A _11186_/S sky130_fd_sc_hd__or2_1
XFILLER_76_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_49_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14728_ _14728_/Q _14728_/CLK _14728_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_60_584 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14659_ hold400/A _14659_/CLK _14659_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07200_ VGND VPWR VPWR VGND _07358_/B _15598_/Q _07230_/S _14387_/Q sky130_fd_sc_hd__mux2_1
X_08180_ VPWR VGND VGND VPWR _08180_/A _08180_/B _08181_/B _08180_/C sky130_fd_sc_hd__nand3_1
X_07131_ VGND VPWR VPWR VGND _09556_/C _09240_/A _09311_/B _08377_/A sky130_fd_sc_hd__or3b_1
X_07964_ VGND VPWR VGND VPWR _07186_/A _07981_/A _07981_/B _07965_/B sky130_fd_sc_hd__o21ba_1
X_13399__516 VPWR VGND VPWR VGND _14674_/CLK clkload9/A sky130_fd_sc_hd__inv_2
XFILLER_56_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07895_ VPWR VGND VPWR VGND _11102_/S _07119_/A clone17/A _07895_/Y sky130_fd_sc_hd__a21oi_1
X_09703_ VGND VPWR VPWR VGND _14340_/D fanout66/X _09710_/S hold662/X sky130_fd_sc_hd__mux2_1
XFILLER_74_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13143__260 VPWR VGND VPWR VGND _14418_/CLK clkload9/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_27_Left_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09634_ VGND VPWR VPWR VGND _14436_/D hold925/X _09637_/S fanout65/X sky130_fd_sc_hd__mux2_1
XFILLER_56_879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09565_ VGND VPWR VPWR VGND _14500_/D hold900/X _09584_/S fanout65/X sky130_fd_sc_hd__mux2_1
X_08516_ VPWR VGND _15328_/D _08516_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
X_09496_ VGND VPWR VPWR VGND _14563_/D fanout61/X _09517_/S hold516/X sky130_fd_sc_hd__mux2_1
X_08447_ VGND VPWR VGND VPWR _15353_/D hold1340/X _08448_/B _08446_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_23_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14026__1143 VPWR VGND VPWR VGND _15398_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_08378_ VPWR VGND VPWR VGND _08378_/Y _08405_/S sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_36_Left_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07329_ _07329_/X _07416_/A _07154_/A _07325_/Y _07966_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_10340_ VPWR VGND VGND VPWR _10340_/X _14385_/Q _12269_/B sky130_fd_sc_hd__or2_1
X_10271_ VGND VPWR VPWR VGND _10271_/X hold586/A _10271_/S hold195/A sky130_fd_sc_hd__mux2_1
X_12010_ VPWR VGND VPWR VGND _12009_/X _12029_/A _12047_/B1 _12010_/X sky130_fd_sc_hd__a21o_1
X_13955__1072 VPWR VGND VPWR VGND _15327_/CLK clkload25/A sky130_fd_sc_hd__inv_2
Xfanout450 VPWR VGND _10737_/C1 _07593_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout461 VPWR VGND VGND VPWR _07592_/Y clone2/A sky130_fd_sc_hd__buf_12
Xfanout472 VGND VPWR _12705_/A2 _12746_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_59_662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Left_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout483 VPWR VGND _12006_/B _12005_/S VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_24_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15700_ VGND VPWR hold151/A uo_out[5] VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout494 VGND VPWR _11965_/S _12191_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_76_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15631_ _15631_/Q clkload49/A _15631_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12843_ VGND VPWR VGND VPWR _12846_/B _15571_/Q _07234_/B _12843_/X sky130_fd_sc_hd__o21ba_1
XFILLER_76_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15562_ _15562_/Q clkload44/A _15562_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12774_ VPWR VGND VGND VPWR _12774_/X _12789_/A _12774_/B sky130_fd_sc_hd__or2_1
X_13192__309 VPWR VGND VPWR VGND _14467_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_13883__1000 VPWR VGND VPWR VGND _15255_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_14513_ hold286/A _14513_/CLK _14513_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15493_ hold844/A _15493_/CLK _15493_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11725_ VGND VPWR VPWR VGND _11725_/X hold703/A _11748_/S hold255/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_54_Left_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14444_ hold520/A _14444_/CLK _14444_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11656_ VGND VPWR VPWR VGND _11656_/X _11653_/X _11948_/S _11652_/X sky130_fd_sc_hd__mux2_1
Xfanout90 VPWR VGND fanout90/X _07600_/X VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_30_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11587_ VGND VPWR VPWR VGND _11587_/X hold851/A _12094_/S hold531/A sky130_fd_sc_hd__mux2_1
X_14375_ hold793/A _14375_/CLK _14375_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10607_ VGND VPWR VPWR VGND _10607_/X _10604_/X _10615_/S _10603_/X sky130_fd_sc_hd__mux2_1
X_10538_ VGND VPWR VPWR VGND _10538_/X hold854/A _10700_/S hold175/A sky130_fd_sc_hd__mux2_1
Xhold909 hold909/X hold909/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13086__203 VPWR VGND VPWR VGND _14329_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_10469_ VGND VPWR VPWR VGND _10470_/B _10468_/Y _10469_/S _10460_/Y sky130_fd_sc_hd__mux2_1
X_12208_ VGND VPWR VPWR VGND _12208_/X hold617/A _12228_/B hold211/A sky130_fd_sc_hd__mux2_1
XFILLER_9_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_9_1027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Left_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12139_ VGND VPWR VPWR VGND _12140_/B _12138_/Y _12139_/S _12130_/Y sky130_fd_sc_hd__mux2_1
X_13127__244 VPWR VGND VPWR VGND _14370_/CLK clkload41/A sky130_fd_sc_hd__inv_2
XFILLER_38_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07680_ VGND VPWR VGND VPWR _07681_/C _07694_/B _07401_/B _07693_/B _07679_/A sky130_fd_sc_hd__a211o_1
XFILLER_52_326 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09350_ VGND VPWR VPWR VGND _09357_/S hold1118/X clone49/X _14696_/D sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_72_Left_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13784__901 VPWR VGND VPWR VGND _15156_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_08301_ VGND VPWR VPWR VGND _09311_/B _09556_/C _09240_/A _09591_/A sky130_fd_sc_hd__or3_2
X_09281_ VGND VPWR VPWR VGND _14760_/D clone49/A _09304_/S hold299/X sky130_fd_sc_hd__mux2_1
X_08232_ VPWR VGND VGND VPWR _08232_/A _08232_/Y _08232_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_1224 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13825__942 VPWR VGND VPWR VGND _15197_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_08163_ VPWR VGND VPWR VGND _08162_/B _08162_/A _08240_/A _08163_/X sky130_fd_sc_hd__a21o_1
X_07114_ VPWR VGND VPWR VGND _09486_/B _15577_/Q sky130_fd_sc_hd__inv_2
X_08094_ VGND VPWR VPWR VGND _08094_/X _08093_/X _08684_/S _07661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08996_ VGND VPWR VGND VPWR _08996_/X _09873_/A _09016_/B1 _15104_/Q _08995_/Y sky130_fd_sc_hd__a211o_1
XFILLER_0_639 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_76_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07947_ VPWR VGND VPWR VGND _15083_/Q _10072_/B _07947_/X _10074_/A0 _07288_/A _07946_/Y
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_802 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1386 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_805 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07878_ VPWR VGND VPWR VGND _07878_/B _07878_/C _07878_/A _07878_/X sky130_fd_sc_hd__or3_1
X_09617_ VGND VPWR VPWR VGND _14451_/D _09825_/A1 _09617_/S hold569/X sky130_fd_sc_hd__mux2_1
X_09548_ VGND VPWR VPWR VGND _14514_/D _09548_/A1 _09555_/S hold194/X sky130_fd_sc_hd__mux2_1
X_09479_ VGND VPWR VPWR VGND _14577_/D _09827_/A1 _09482_/S hold349/X sky130_fd_sc_hd__mux2_1
X_11510_ VGND VPWR VPWR VGND _15087_/D _11509_/X _11538_/S _15087_/Q sky130_fd_sc_hd__mux2_1
XFILLER_12_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12490_ VPWR VGND _12490_/X _12489_/X _12485_/X _12472_/S _12481_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11441_ VGND VPWR VGND VPWR _11440_/Y _11340_/A _11441_/Y _12845_/B sky130_fd_sc_hd__a21oi_4
X_11372_ VGND VPWR VPWR VGND _11372_/X _11371_/X _11387_/S _14845_/Q sky130_fd_sc_hd__mux2_1
X_13568__685 VPWR VGND VPWR VGND _14899_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_14160_ hold395/A _14160_/CLK _14160_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10323_ VPWR VGND VPWR VGND _10322_/X _10851_/A _11263_/C1 _10323_/X sky130_fd_sc_hd__a21o_1
X_10254_ VGND VPWR VPWR VGND _10254_/X _14351_/Q _10924_/B hold675/A sky130_fd_sc_hd__mux2_1
XFILLER_59_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10185_ VPWR VGND VGND VPWR _10185_/X _10703_/A _10185_/B sky130_fd_sc_hd__or2_1
X_12960__77 VPWR VGND VPWR VGND _14203_/CLK clkload21/A sky130_fd_sc_hd__inv_2
Xfanout280 VGND VPWR fanout282/X _11262_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_43_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14993_ hold332/A _14993_/CLK _14993_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_3_Left_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout291 VPWR VGND _10521_/B _10520_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_15614_ _15614_/Q clkload27/A _15614_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12826_ VPWR VGND VGND VPWR _12831_/A _12826_/B _12826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15545_ _15545_/Q clkload32/A _15545_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12757_ VGND VPWR VGND VPWR _15546_/D _10060_/A _15546_/Q _09976_/B _12756_/Y sky130_fd_sc_hd__o211a_1
X_13809__926 VPWR VGND VPWR VGND _15181_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_12688_ VGND VPWR VPWR VGND _12688_/X _14217_/Q _12689_/S hold222/A sky130_fd_sc_hd__mux2_1
X_15476_ _15476_/Q clkload33/A _15476_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11708_ VGND VPWR VGND VPWR _11708_/X _11705_/X _11707_/X _12489_/A1 _12485_/C1 sky130_fd_sc_hd__a211o_1
X_14427_ hold998/A _14427_/CLK _14427_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11639_ VPWR VGND _11639_/X _11638_/X _11634_/X _12102_/S _11630_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14358_ hold875/A _14358_/CLK _14358_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold706 hold706/X hold706/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 hold717/X hold717/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 hold728/X hold728/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ hold152/A _14289_/CLK _14289_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold739 hold739/X hold739/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08850_ VGND VPWR VPWR VGND _15163_/D fanout96/X _08850_/S hold626/X sky130_fd_sc_hd__mux2_1
X_07801_ _07915_/B _07722_/Y _07800_/A _07800_/B _07938_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xhold1406 hold1406/X _15096_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13361__478 VPWR VGND VPWR VGND _14636_/CLK clkload8/A sky130_fd_sc_hd__inv_2
Xhold1439 hold1439/X hold837/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 hold1428/X hold988/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14025__1142 VPWR VGND VPWR VGND _15397_/CLK clkload54/A sky130_fd_sc_hd__inv_2
Xhold1417 hold1417/X _15079_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08781_ VPWR VGND VPWR VGND _08781_/Y _08811_/S sky130_fd_sc_hd__inv_2
X_07732_ VPWR VGND VGND VPWR _15557_/Q _07998_/B _07734_/B sky130_fd_sc_hd__nand2_1
X_07663_ VGND VPWR _07664_/B _07663_/B _07663_/A _07665_/A VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_53_657 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09402_ VGND VPWR VPWR VGND _14647_/D hold472/X _09414_/S fanout15/X sky130_fd_sc_hd__mux2_1
XFILLER_20_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07594_ VGND VPWR VPWR VGND _08151_/B _08073_/B _10728_/S _07591_/A sky130_fd_sc_hd__mux2_4
X_09333_ VGND VPWR VPWR VGND _14711_/D hold502/X _09345_/S fanout17/X sky130_fd_sc_hd__mux2_1
X_13954__1071 VPWR VGND VPWR VGND _15326_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_09264_ VGND VPWR VPWR VGND _14779_/D fanout12/X _09275_/S hold601/X sky130_fd_sc_hd__mux2_1
X_13255__372 VPWR VGND VPWR VGND _14530_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_08215_ VPWR VGND VPWR VGND _08174_/Y _15336_/Q _08491_/A _08215_/X _14839_/Q sky130_fd_sc_hd__a22o_1
X_09195_ VGND VPWR VPWR VGND _14896_/D hold649/X _09197_/S _09229_/A0 sky130_fd_sc_hd__mux2_1
X_08146_ VGND VPWR _08146_/B _12772_/A _08146_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_08077_ VPWR VGND _08078_/B _08145_/A _15552_/Q _15553_/Q _15554_/Q VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_49_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13602__719 VPWR VGND VPWR VGND _14942_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
XFILLER_1_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_1448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08979_ VGND VPWR VGND VPWR _15111_/D hold1044/X _08985_/A2 _08978_/X _08955_/A sky130_fd_sc_hd__o211a_1
XFILLER_29_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11990_ VPWR VGND VPWR VGND _11989_/X _12008_/C1 _11988_/X _11990_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_687 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10941_ VPWR VGND VPWR VGND _10940_/X _11181_/A1 _10939_/X _10941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_32 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10872_ VPWR VGND VGND VPWR _10872_/X _14304_/Q _11241_/S sky130_fd_sc_hd__or2_1
X_12611_ VPWR VGND VPWR VGND _12610_/X _12740_/A1 _12609_/X _12611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15330_ _15330_/Q _15330_/CLK _15330_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12542_ VPWR VGND VGND VPWR _12542_/X _12665_/S _12542_/B sky130_fd_sc_hd__or2_1
X_15261_ _15698_/A _15261_/CLK _15261_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12473_ VPWR VGND VGND VPWR _12473_/A _12473_/B _12473_/Y sky130_fd_sc_hd__nor2_1
X_11424_ VGND VPWR VGND VPWR _11424_/X _14927_/Q _11303_/A _11431_/A2 sky130_fd_sc_hd__a21bo_1
X_14212_ _14212_/Q _14212_/CLK _14212_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_8 _08059_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15192_ hold510/A _15192_/CLK _15192_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14143_ hold714/A _14143_/CLK hold715/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11355_ VGND VPWR VPWR VGND _11355_/X _14933_/Q _11355_/S hold1297/X sky130_fd_sc_hd__mux2_1
XFILLER_10_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10306_ VGND VPWR VPWR VGND _10306_/X hold912/A _11098_/S hold551/A sky130_fd_sc_hd__mux2_1
X_11286_ VPWR VGND _14811_/D _11286_/B _11382_/S VPWR VGND sky130_fd_sc_hd__and2_1
X_10237_ VGND VPWR VPWR VGND _10237_/X _10234_/X _10911_/S _10233_/X sky130_fd_sc_hd__mux2_1
X_10168_ VGND VPWR VPWR VGND _10168_/X hold666/A _10169_/B hold257/A sky130_fd_sc_hd__mux2_1
XFILLER_0_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13198__315 VPWR VGND VPWR VGND _14473_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_10099_ VGND VPWR VPWR VGND _10100_/B _10098_/Y _10617_/S _10090_/Y sky130_fd_sc_hd__mux2_1
X_14976_ hold678/A _14976_/CLK _14976_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13239__356 VPWR VGND VPWR VGND _14514_/CLK clkload10/A sky130_fd_sc_hd__inv_2
XFILLER_62_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12809_ VPWR VGND VGND VPWR _12809_/X _12817_/A _12809_/B sky130_fd_sc_hd__or2_1
XFILLER_31_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15528_ hold166/A _15528_/CLK _15528_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1087 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08000_ VGND VPWR _08023_/A _08000_/Y _15558_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_15459_ VGND VPWR VGND VPWR _15459_/Q _15459_/D clkload10/A sky130_fd_sc_hd__dfxtp_4
Xhold536 hold536/X hold536/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 hold514/X hold514/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 hold503/X hold503/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 hold525/X hold525/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ VGND VPWR _09954_/C _09951_/Y _14127_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold569 hold569/X hold569/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 hold547/X hold547/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 hold558/X hold558/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ VPWR VGND VGND VPWR _08902_/A _08902_/Y _08902_/B sky130_fd_sc_hd__nand2_1
X_09882_ VPWR VGND VGND VPWR _09882_/A _09882_/B _14149_/D sky130_fd_sc_hd__nor2_1
Xhold1225 _14836_/D _11349_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 hold1214/X _14279_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1203 hold1203/X _14440_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08833_ VGND VPWR VPWR VGND _15180_/D fanout37/X _08842_/S hold646/X sky130_fd_sc_hd__mux2_1
Xhold1247 hold1247/X _14956_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 _15160_/D _08865_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1236 hold1236/X _15358_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ VGND VPWR VPWR VGND _15242_/D fanout29/X _08772_/S hold273/X sky130_fd_sc_hd__mux2_1
X_07715_ VPWR VGND VPWR VGND _07827_/D _15589_/Q _07714_/X _07717_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_900 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1269 hold1269/X _14963_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08695_ VGND VPWR VGND VPWR _15283_/D hold953/X _08701_/A2 _08694_/X _11937_/C1 sky130_fd_sc_hd__o211a_1
X_07646_ VGND VPWR VGND VPWR _07914_/B1 _07659_/B _07645_/X _07418_/B sky130_fd_sc_hd__o21ba_4
X_07577_ VPWR VGND VGND VPWR _07577_/A _07578_/B _07577_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_1105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09316_ VGND VPWR VPWR VGND _09327_/S hold1099/X fanout81/X _14728_/D sky130_fd_sc_hd__mux2_2
X_09247_ VGND VPWR VPWR VGND _14796_/D _09269_/S fanout76/X hold1223/X sky130_fd_sc_hd__mux2_4
X_09178_ VGND VPWR VPWR VGND _14913_/D hold585/X _09194_/S clone6/A sky130_fd_sc_hd__mux2_1
X_13032__149 VPWR VGND VPWR VGND _14275_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_08129_ VGND VPWR VPWR VGND _15522_/D fanout5/X _08300_/S hold191/X sky130_fd_sc_hd__mux2_1
X_11140_ VGND VPWR VGND VPWR _11140_/X _11139_/X _11138_/X _11189_/A1 _11254_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_27_1212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11071_ VGND VPWR VPWR VGND _11071_/X hold698/A _11186_/S hold306/A sky130_fd_sc_hd__mux2_1
X_12930__47 VPWR VGND VPWR VGND _14173_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_10022_ VPWR VGND VGND VPWR _10024_/C _10022_/B _15624_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14830_ _14830_/Q _14832_/CLK _14830_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11973_ VPWR VGND VGND VPWR _11973_/A _11973_/Y _11973_/B sky130_fd_sc_hd__nand2_1
X_14761_ hold249/A _14761_/CLK _14761_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_17_646 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14692_ hold469/A _14692_/CLK _14692_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10924_ VPWR VGND VGND VPWR _10924_/X hold168/A _10924_/B sky130_fd_sc_hd__or2_1
X_13730__847 VPWR VGND VPWR VGND _15102_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_10855_ VPWR VGND VGND VPWR _10852_/X _10854_/X _11209_/S _10855_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15313_ hold905/A _15313_/CLK _15313_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10786_ VGND VPWR VPWR VGND _10786_/X _14622_/Q _11216_/S _14654_/Q sky130_fd_sc_hd__mux2_1
XFILLER_40_671 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12525_ VGND VPWR VGND VPWR _12525_/X _15024_/Q _12743_/A2 _12735_/S _12524_/X sky130_fd_sc_hd__o211a_1
X_13583__700 VPWR VGND VPWR VGND _14914_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_14024__1141 VPWR VGND VPWR VGND _15396_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_15244_ hold258/A _15244_/CLK _15244_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12456_ VGND VPWR VPWR VGND _12460_/B hold623/A _12477_/B hold400/A sky130_fd_sc_hd__mux2_1
X_11407_ VPWR VGND VGND VPWR _14856_/Q _11410_/B _14855_/Q sky130_fd_sc_hd__nand2_1
X_15175_ hold417/A _15175_/CLK _15175_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12387_ VGND VPWR VGND VPWR _12387_/X _12720_/A1 _12383_/X _12386_/X _12720_/C1 sky130_fd_sc_hd__o211a_1
X_11338_ VGND VPWR _11338_/B _11338_/Y _14832_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_14126_ _14126_/Q _14126_/CLK _14126_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13624__741 VPWR VGND VPWR VGND _14964_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_11269_ VPWR VGND VGND VPWR _11545_/B _15432_/Q _11269_/B sky130_fd_sc_hd__or2_1
X_13953__1070 VPWR VGND VPWR VGND _15325_/CLK clkload26/A sky130_fd_sc_hd__inv_2
XFILLER_55_708 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_11_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_782 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_36_900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07500_ VPWR VGND VGND VPWR _07551_/A _07500_/Y _07551_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14959_ hold729/A _14959_/CLK _14959_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08480_ VPWR VGND VGND VPWR _08480_/X _15336_/Q _08482_/B sky130_fd_sc_hd__or2_1
X_07431_ VPWR VGND _07433_/A _07511_/B _15461_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_56_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07362_ VPWR VGND VPWR VGND _08275_/A _08258_/B _10061_/A _07362_/Y sky130_fd_sc_hd__a21oi_1
X_09101_ VGND VPWR VPWR VGND _14994_/D _09122_/S hold1106/X fanout72/X sky130_fd_sc_hd__mux2_4
X_07293_ VGND VPWR VGND VPWR _07291_/X _07820_/A _07293_/B sky130_fd_sc_hd__nand2b_2
X_09032_ VGND VPWR VPWR VGND _15058_/D _09053_/S hold1121/X fanout72/X sky130_fd_sc_hd__mux2_4
Xhold311 hold311/X hold311/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold300 hold300/X hold300/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 hold333/X hold333/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 hold344/X hold344/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13367__484 VPWR VGND VPWR VGND _14642_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
Xhold322 hold322/X hold322/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold355 hold355/X hold355/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 hold377/X hold377/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 hold366/X hold366/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout824 VGND VPWR _08571_/B fanout824/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout802 VPWR VGND fanout802/X _14765_/Q VPWR VGND sky130_fd_sc_hd__buf_2
X_09934_ VPWR VGND VPWR VGND _09919_/Y _08498_/Y hold239/X _09934_/Y sky130_fd_sc_hd__a21oi_1
Xhold399 hold399/X hold399/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 VPWR VGND VPWR VGND _08717_/C1 _12159_/C1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold388 hold388/X hold388/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout835 VPWR VGND VPWR VGND _09017_/A _09976_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09865_ VGND VPWR VPWR VGND _14157_/D hold636/X _09865_/S _09865_/A0 sky130_fd_sc_hd__mux2_1
Xfanout857 VGND VPWR _07327_/X _08182_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold1000 hold1000/X _15268_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout846 VGND VPWR _07422_/X _08293_/A3 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold1011 hold1011/X _15121_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 VPWR VGND _07507_/B _07511_/B VPWR VGND sky130_fd_sc_hd__buf_2
Xhold1022 hold1022/X _15001_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ VPWR VGND VGND VPWR _09095_/B _08816_/Y _09694_/A sky130_fd_sc_hd__nor2_2
Xfanout879 VPWR VGND VPWR VGND _12855_/A0 _15579_/Q sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1033 hold1033/X _15005_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1044 hold1044/X _15111_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ VGND VPWR VPWR VGND _14253_/D _09865_/A0 _09798_/S hold1040/X sky130_fd_sc_hd__mux2_1
Xhold1055 hold1055/X _15019_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 hold1066/X _15007_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 hold1077/X _15503_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 hold1099/X _14728_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 hold1088/X _15027_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ VPWR VGND VGND VPWR _08747_/X _08747_/A _08776_/S sky130_fd_sc_hd__or2_1
X_08678_ VGND VPWR VPWR VGND _08678_/X _14399_/Q _08684_/S _14383_/Q sky130_fd_sc_hd__mux2_1
XFILLER_27_977 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07629_ VPWR VGND VPWR VGND _07629_/B _07629_/C _07629_/A clone45/A sky130_fd_sc_hd__or3_4
X_10640_ VGND VPWR VPWR VGND _10640_/X hold700/A _10720_/S hold273/A sky130_fd_sc_hd__mux2_1
XFILLER_42_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10571_ VPWR VGND VPWR VGND _10570_/X _10745_/C1 _10569_/X _10571_/Y sky130_fd_sc_hd__a21oi_1
X_12310_ VGND VPWR VPWR VGND _12310_/X hold829/A _12318_/S hold317/A sky130_fd_sc_hd__mux2_1
X_12241_ VGND VPWR VGND VPWR _12241_/X _12240_/X _12239_/X _12581_/S _12702_/C1 sky130_fd_sc_hd__a211o_1
X_13608__725 VPWR VGND VPWR VGND _14948_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_12172_ VPWR VGND VGND VPWR _12172_/X _12174_/S _12172_/B sky130_fd_sc_hd__or2_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11123_ VPWR VGND VGND VPWR _11123_/X _11143_/S _11123_/B sky130_fd_sc_hd__or2_1
X_11054_ VGND VPWR VPWR VGND _11054_/X hold575/A _11054_/S hold373/A sky130_fd_sc_hd__mux2_1
X_10005_ VPWR VGND VGND VPWR _10007_/B _10005_/B _15617_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14813_ _14813_/Q clkload20/A _14813_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13160__277 VPWR VGND VPWR VGND _14435_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_11956_ VGND VPWR VPWR VGND _11956_/X hold830/A _11964_/S hold356/A sky130_fd_sc_hd__mux2_1
X_14744_ hold444/A _14744_/CLK _14744_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10907_ VGND VPWR VPWR VGND _10907_/X _14209_/Q _10919_/S _15217_/Q sky130_fd_sc_hd__mux2_1
XFILLER_60_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14675_ hold686/A _14675_/CLK _14675_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11887_ VPWR VGND VPWR VGND _11886_/X _12175_/A1 _11885_/X _11887_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_1160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10838_ VGND VPWR VGND VPWR _10838_/X _11104_/B1 _10833_/X _10837_/X _11209_/S sky130_fd_sc_hd__o211a_1
X_10769_ VGND VPWR VPWR VGND _10769_/X _10768_/X _11092_/S _10767_/X sky130_fd_sc_hd__mux2_1
X_12508_ VPWR VGND VPWR VGND _12507_/X _12666_/A1 _12506_/X _12508_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13054__171 VPWR VGND VPWR VGND _14297_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_15227_ hold160/A _15227_/CLK _15227_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12439_ VGND VPWR VPWR VGND _12439_/X _12438_/X _12655_/S _12437_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_1344 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_59_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15158_ _15158_/Q _15158_/CLK _15158_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12892__9 VPWR VGND VPWR VGND _14134_/CLK clkload25/A sky130_fd_sc_hd__inv_2
Xfanout109 VGND VPWR _08266_/X _09865_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07980_ VPWR VGND VPWR VGND _12375_/S _08286_/A _07598_/Y _07994_/A sky130_fd_sc_hd__a21oi_1
X_15089_ _15089_/Q clkload36/A _15089_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09650_ VGND VPWR VPWR VGND _14420_/D hold885/X _09657_/S fanout5/X sky130_fd_sc_hd__mux2_1
X_13401__518 VPWR VGND VPWR VGND _14676_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_08601_ VGND VPWR VGND VPWR _08601_/X _08605_/A _08615_/B1 hold1052/X _08600_/Y sky130_fd_sc_hd__a211o_1
X_09581_ VGND VPWR VPWR VGND _14484_/D hold1030/X _09588_/S fanout6/X sky130_fd_sc_hd__mux2_1
X_08532_ VPWR VGND VPWR VGND _08534_/B1 _15319_/Q _08540_/A2 _08533_/B hold1436/X
+ sky130_fd_sc_hd__a22o_1
X_08463_ VGND VPWR VGND VPWR _15345_/D hold1176/X _08483_/A2 _08462_/X _11974_/C1
+ sky130_fd_sc_hd__o211a_1
X_07414_ VPWR VGND VGND VPWR _08198_/S _07414_/Y _10072_/A sky130_fd_sc_hd__nor2_2
X_08394_ VGND VPWR VPWR VGND _15383_/D fanout37/X _08409_/S hold633/X sky130_fd_sc_hd__mux2_1
X_07345_ VGND VPWR _07345_/X _07971_/A _15461_/Q _07345_/C VPWR VGND sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_30_clk _14832_/CLK clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07276_ VPWR VGND VPWR VGND _07186_/A _07181_/Y _07182_/A _07916_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_1400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09015_ VGND VPWR VGND VPWR _15099_/D hold1057/X _09015_/A2 _09014_/X _11327_/A sky130_fd_sc_hd__o211a_1
Xhold152 hold152/X hold152/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_619 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold163 hold163/X hold163/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/X hold185/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/X hold174/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ VPWR VGND VGND VPWR _09917_/A _09917_/B _14138_/D sky130_fd_sc_hd__nor2_1
Xfanout621 VPWR VGND _09861_/S _09864_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xhold196 hold196/X hold196/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout632 VPWR VGND _09684_/S _09660_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout610 VGND VPWR _08251_/S _08267_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_12900__17 VPWR VGND VPWR VGND _14142_/CLK clkload29/A sky130_fd_sc_hd__inv_2
Xfanout676 VPWR VGND _09122_/S _09125_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout643 _09587_/S _09557_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout665 _09231_/S _09229_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout654 VPWR VGND _09478_/S _09451_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout698 VPWR VGND _08918_/B _08868_/B VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout687 VPWR VGND _08338_/S _08330_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09848_ VGND VPWR VPWR VGND _14174_/D _09864_/S hold1163/X clone44/X sky130_fd_sc_hd__mux2_4
XFILLER_37_22 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09779_ VGND VPWR VPWR VGND _14270_/D clone6/X _09795_/S hold790/X sky130_fd_sc_hd__mux2_1
X_14023__1140 VPWR VGND VPWR VGND _15395_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_11810_ VGND VPWR VPWR VGND _11810_/X _11809_/X _11810_/S _11808_/X sky130_fd_sc_hd__mux2_1
X_12790_ VPWR VGND VGND VPWR _12790_/A _12790_/Y _12790_/B sky130_fd_sc_hd__nand2_1
X_11741_ VGND VPWR VGND VPWR _11741_/X _12415_/C1 _11736_/X _11740_/X _12864_/A1 sky130_fd_sc_hd__o211a_1
X_11672_ VGND VPWR VPWR VGND _11672_/X hold984/A _11965_/S hold653/A sky130_fd_sc_hd__mux2_1
X_14460_ hold617/A _14460_/CLK _14460_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13038__155 VPWR VGND VPWR VGND _14281_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_14391_ _14391_/Q clkload13/A _14391_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10623_ VGND VPWR VPWR VGND _10623_/X hold800/A _10632_/B hold440/A sky130_fd_sc_hd__mux2_1
XFILLER_23_980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_clk clkload28/A clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_10554_ VGND VPWR VPWR VGND _10557_/B hold844/A _10554_/S hold546/A sky130_fd_sc_hd__mux2_1
X_13842__959 VPWR VGND VPWR VGND _15214_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_10485_ VGND VPWR VGND VPWR _10485_/X _15009_/Q _10688_/A2 _10484_/X _10677_/S sky130_fd_sc_hd__o211a_1
X_15012_ _15012_/Q _15012_/CLK _15012_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12224_ VPWR VGND VGND VPWR _12224_/X hold316/A _12227_/S sky130_fd_sc_hd__or2_1
X_12155_ VGND VPWR VPWR VGND _12155_/X hold756/A _12155_/S hold166/A sky130_fd_sc_hd__mux2_1
X_11106_ VGND VPWR VPWR VGND _11110_/B hold691/A _11109_/S _15058_/Q sky130_fd_sc_hd__mux2_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13695__812 VPWR VGND VPWR VGND _15035_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_42_1304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12086_ VGND VPWR VPWR VGND _12090_/B hold521/A _12086_/S hold667/A sky130_fd_sc_hd__mux2_1
X_11037_ VGND VPWR VGND VPWR _11037_/X _11034_/X _11036_/X _11252_/C1 _11245_/A1 sky130_fd_sc_hd__a211o_1
X_13736__853 VPWR VGND VPWR VGND _15108_/CLK clkload46/A sky130_fd_sc_hd__inv_2
XFILLER_75_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11939_ VPWR VGND VGND VPWR _11939_/X hold545/A _11950_/B sky130_fd_sc_hd__or2_1
X_14119__1236 VPWR VGND VPWR VGND _15538_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_14727_ hold598/A _14727_/CLK _14727_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_33_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14658_ hold559/A _14658_/CLK _14658_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07130_ VPWR VGND VPWR VGND _09486_/B _09198_/B _09164_/A _09799_/A sky130_fd_sc_hd__or3_4
X_14589_ hold256/A _14589_/CLK _14589_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clkload21/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12966__83 VPWR VGND VPWR VGND _14209_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_60_1415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07963_ VPWR VGND VPWR VGND _07962_/Y _12833_/A _07960_/X _07963_/X sky130_fd_sc_hd__a21o_1
X_07894_ VGND VPWR VGND VPWR _07894_/X clone18/A _15141_/Q _07892_/Y sky130_fd_sc_hd__a21bo_1
X_09702_ VGND VPWR VPWR VGND _14341_/D fanout69/X _09710_/S hold946/X sky130_fd_sc_hd__mux2_1
X_09633_ VGND VPWR VPWR VGND _14437_/D hold1037/X _09637_/S fanout71/X sky130_fd_sc_hd__mux2_1
X_13479__596 VPWR VGND VPWR VGND _14754_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_09564_ VGND VPWR VPWR VGND _14501_/D hold1045/X _09584_/S fanout69/X sky130_fd_sc_hd__mux2_1
X_08515_ VPWR VGND VPWR VGND _08534_/B1 _15327_/Q _08503_/A _08516_/B hold1421/X sky130_fd_sc_hd__a22o_1
XFILLER_58_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_51_530 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09495_ VGND VPWR VPWR VGND _14564_/D fanout66/X _09514_/S hold740/X sky130_fd_sc_hd__mux2_1
X_08446_ VPWR VGND VGND VPWR _08446_/X _15353_/Q _08488_/B sky130_fd_sc_hd__or2_1
X_08377_ VPWR VGND VGND VPWR _09694_/A _08377_/Y _08377_/A sky130_fd_sc_hd__nor2_2
XFILLER_11_416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07328_ VPWR VGND VGND VPWR _07328_/Y _11535_/A _07328_/B sky130_fd_sc_hd__nand2_2
XFILLER_20_950 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13932__1049 VPWR VGND VPWR VGND _15304_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_07259_ VPWR VGND VPWR VGND _07260_/B _07271_/B sky130_fd_sc_hd__inv_2
X_10270_ VGND VPWR VPWR VGND _10270_/X hold689/A _10602_/S hold221/A sky130_fd_sc_hd__mux2_1
Xfanout440 VGND VPWR _11023_/A1 _11096_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13423__540 VPWR VGND VPWR VGND _14698_/CLK clkload38/A sky130_fd_sc_hd__inv_2
Xfanout451 VPWR VGND _11255_/C1 _12869_/A1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout473 VGND VPWR _12080_/A2 _12705_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout484 VGND VPWR _12005_/S _12117_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout462 VGND VPWR _12040_/A2 _12188_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout495 VGND VPWR _11965_/S _12190_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_15630_ _15630_/Q clkload49/A _15630_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_73_154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12842_ VPWR VGND _12842_/X _12842_/B _15570_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_15561_ _15561_/Q clkload44/A _15561_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12773_ VGND VPWR VGND VPWR _12773_/X _12788_/S _12772_/Y _08145_/Y _12790_/A sky130_fd_sc_hd__a211o_1
XFILLER_55_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11724_ VGND VPWR VPWR VGND _11728_/B hold753/A _11748_/S hold347/A sky130_fd_sc_hd__mux2_1
X_15492_ hold669/A _15492_/CLK _15492_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14512_ hold203/A _14512_/CLK _14512_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11655_ VGND VPWR VGND VPWR _11655_/X _11968_/S _11651_/X _11654_/X _12189_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_42_596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14443_ hold789/A _14443_/CLK _14443_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13272__389 VPWR VGND VPWR VGND _14547_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
Xfanout91 VPWR VGND fanout91/X fanout92/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout80 VGND VPWR clone45/A fanout80/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_14374_ _14374_/Q _14374_/CLK _14374_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11586_ VGND VPWR VPWR VGND _11586_/X hold878/A _11998_/S hold464/A sky130_fd_sc_hd__mux2_1
X_10606_ VGND VPWR VGND VPWR _10606_/X _10614_/A1 _10602_/X _10605_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
X_10537_ VGND VPWR VPWR VGND _10537_/X _10536_/X _10703_/A _10535_/X sky130_fd_sc_hd__mux2_1
X_10468_ VPWR VGND VPWR VGND _10467_/X _10706_/C1 _10466_/X _10468_/Y sky130_fd_sc_hd__a21oi_1
X_12207_ VGND VPWR VPWR VGND _12207_/X _14204_/Q _12228_/B hold550/A sky130_fd_sc_hd__mux2_1
X_10399_ VGND VPWR VPWR VGND _10399_/X _10398_/X _10677_/S _10397_/X sky130_fd_sc_hd__mux2_1
X_13166__283 VPWR VGND VPWR VGND _14441_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_12138_ VPWR VGND VPWR VGND _12137_/X _12212_/A1 _12136_/X _12138_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_670 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_78_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12069_ VGND VPWR VPWR VGND _12069_/X _12068_/X _12069_/S _12067_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_1_clk clkload6/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_38_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_688 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09280_ VGND VPWR VPWR VGND _14761_/D fanout85/X _09304_/S hold249/X sky130_fd_sc_hd__mux2_1
X_08300_ VGND VPWR VPWR VGND _15513_/D fanout96/X _08300_/S hold192/X sky130_fd_sc_hd__mux2_1
X_08231_ VGND VPWR VPWR VGND _15517_/D _09689_/A0 _08231_/S hold511/X sky130_fd_sc_hd__mux2_1
X_08162_ VPWR VGND VGND VPWR _08162_/A _08162_/B _08162_/Y sky130_fd_sc_hd__nor2_1
X_13864__981 VPWR VGND VPWR VGND _15236_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_08093_ VPWR VGND VPWR VGND _08252_/A2 _15342_/Q _08253_/A2 _08093_/X _15147_/Q sky130_fd_sc_hd__a22o_1
X_07113_ VPWR VGND VPWR VGND _07113_/Y _15591_/Q sky130_fd_sc_hd__inv_2
Xclkload50 clkload50/Y clkload50/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
X_13407__524 VPWR VGND VPWR VGND _14682_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_08995_ VPWR VGND VGND VPWR _09890_/A _08995_/B _08995_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07946_ VPWR VGND VGND VPWR _07946_/A _07972_/B _07946_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07877_ VGND VPWR VGND VPWR _07878_/C _07087_/Y _07306_/B _07900_/A _07817_/A sky130_fd_sc_hd__o211a_1
X_09616_ VGND VPWR VPWR VGND _14452_/D fanout7/A _09617_/S hold538/X sky130_fd_sc_hd__mux2_1
X_09547_ VGND VPWR VPWR VGND _14515_/D _09547_/A1 _09553_/S hold381/X sky130_fd_sc_hd__mux2_1
X_09478_ VGND VPWR VPWR VGND _14578_/D _09860_/A0 _09478_/S hold173/X sky130_fd_sc_hd__mux2_1
X_08429_ VGND VPWR VGND VPWR _15362_/D hold728/X _08485_/A2 _08428_/X _11388_/S sky130_fd_sc_hd__o211a_1
XFILLER_51_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_50_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11440_ VPWR VGND VGND VPWR _15640_/Q _11440_/Y _11440_/B sky130_fd_sc_hd__nand2_1
Xclkload0 clkload0/X clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_11371_ VGND VPWR VPWR VGND _11371_/X _14844_/Q _11392_/B _14812_/Q sky130_fd_sc_hd__mux2_1
X_10322_ VGND VPWR VPWR VGND _10322_/X hold859/A _11261_/B hold491/A sky130_fd_sc_hd__mux2_1
X_10253_ VGND VPWR VPWR VGND _10253_/X hold839/A _10924_/B hold638/A sky130_fd_sc_hd__mux2_1
X_14118__1235 VPWR VGND VPWR VGND _15537_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_10184_ VGND VPWR VPWR VGND _10184_/X hold426/A _10479_/S hold355/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout270 VPWR VGND _12473_/A _07912_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout281 VPWR VGND _11215_/A2 fanout282/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout292 VPWR VGND _10632_/B _10520_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_14992_ hold358/A _14992_/CLK _14992_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_62_614 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13200__317 VPWR VGND VPWR VGND _14475_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XFILLER_76_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12825_ VGND VPWR VPWR VGND _12825_/X _07886_/B _12829_/S _07889_/B sky130_fd_sc_hd__mux2_1
X_15613_ _15613_/Q clkload27/A _15613_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15544_ _15544_/Q _15544_/CLK _15544_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12756_ VGND VPWR _12829_/S _12755_/X _12756_/Y _08247_/X VPWR VGND sky130_fd_sc_hd__o21ai_1
X_12687_ VGND VPWR VPWR VGND _12687_/X hold557/A _12689_/S hold323/A sky130_fd_sc_hd__mux2_1
X_15475_ _15475_/Q clkload39/A _15475_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_13848__965 VPWR VGND VPWR VGND _15220_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_11707_ VGND VPWR VGND VPWR _11707_/X hold997/A _12488_/A2 _12470_/S _11706_/X sky130_fd_sc_hd__o211a_1
X_11638_ VGND VPWR VGND VPWR _11638_/X _11635_/X _11637_/X _11638_/A1 _12101_/A1 sky130_fd_sc_hd__a211o_1
X_14426_ hold874/A _14426_/CLK _14426_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14357_ hold929/A _14357_/CLK _14357_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold707 hold707/X hold707/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 hold718/X hold718/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14002__1119 VPWR VGND VPWR VGND _15374_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_11569_ VGND VPWR VPWR VGND _11569_/X hold897/A _12094_/S hold625/A sky130_fd_sc_hd__mux2_1
X_12936__53 VPWR VGND VPWR VGND _14179_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_14288_ hold240/A _14288_/CLK _14288_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold729 hold729/X hold729/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_41_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1407 hold1407/X _14927_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08780_ VPWR VGND VGND VPWR _09591_/A _08780_/Y _09799_/A sky130_fd_sc_hd__nor2_2
X_07800_ VPWR VGND VGND VPWR _07939_/A _07800_/A _07800_/B sky130_fd_sc_hd__or2_1
Xhold1418 hold1418/X _15327_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 _08955_/B _08954_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07731_ VPWR VGND VPWR VGND _07827_/D _15584_/Q _07714_/X _07734_/B sky130_fd_sc_hd__a21o_1
X_13931__1048 VPWR VGND VPWR VGND _15303_/CLK clkload30/A sky130_fd_sc_hd__inv_2
XFILLER_65_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07662_ VGND VPWR VGND VPWR clone17/X _07418_/B _07661_/X _07673_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07593_ VGND VPWR VGND VPWR _07593_/X _15144_/Q _15355_/Q _08495_/A2 clone18/X sky130_fd_sc_hd__a22o_4
XFILLER_0_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09401_ VGND VPWR VPWR VGND _14648_/D hold654/X _09406_/S fanout19/X sky130_fd_sc_hd__mux2_1
XFILLER_53_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09332_ VGND VPWR VPWR VGND _14712_/D hold634/X _09336_/S fanout21/X sky130_fd_sc_hd__mux2_1
X_09263_ VGND VPWR VPWR VGND _14780_/D fanout16/X _09275_/S hold854/X sky130_fd_sc_hd__mux2_1
XFILLER_33_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08214_ VPWR VGND VGND VPWR _08214_/X _08214_/A _08214_/B sky130_fd_sc_hd__or2_1
X_09194_ VGND VPWR VPWR VGND _14897_/D hold499/X _09194_/S _09228_/A0 sky130_fd_sc_hd__mux2_1
X_08145_ VPWR VGND VGND VPWR _08145_/A _08145_/B _08145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08076_ VGND VPWR _08076_/B _08076_/Y _08076_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13641__758 VPWR VGND VPWR VGND _14981_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_66_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08978_ VGND VPWR VGND VPWR _08978_/X _15478_/Q _08972_/A hold954/X _08977_/Y sky130_fd_sc_hd__a211o_1
XFILLER_60_1020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_1370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07929_ VPWR VGND VPWR VGND _08002_/B1 _15625_/Q _07929_/A2 _07933_/A _15589_/Q sky130_fd_sc_hd__a22o_1
X_13494__611 VPWR VGND VPWR VGND _14769_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_5_1278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10940_ VGND VPWR VPWR VGND _10940_/X _10937_/X _11170_/S _10936_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10871_ VGND VPWR VPWR VGND _10871_/X _14789_/Q _10885_/S _14240_/Q sky130_fd_sc_hd__mux2_1
XFILLER_32_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12610_ VGND VPWR VPWR VGND _12610_/X _12607_/X _12624_/S _12606_/X sky130_fd_sc_hd__mux2_1
X_13535__652 VPWR VGND VPWR VGND _14866_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XFILLER_73_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12541_ VGND VPWR VPWR VGND _12541_/X hold658/A _12652_/S hold296/A sky130_fd_sc_hd__mux2_1
X_15260_ _15260_/Q _15260_/CLK _15260_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12472_ VGND VPWR VPWR VGND _12473_/B _12471_/Y _12472_/S _12463_/Y sky130_fd_sc_hd__mux2_1
X_11423_ VGND VPWR VGND VPWR _14926_/D hold1407/X _11431_/A2 _11422_/X _11431_/C1
+ sky130_fd_sc_hd__o211a_1
X_14211_ _14211_/Q _14211_/CLK _14211_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_9 _07978_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_15191_ hold537/A _15191_/CLK _15191_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14142_ _14142_/Q _14142_/CLK _14142_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11354_ VGND VPWR VPWR VGND _11354_/X _14932_/Q _11355_/S hold1255/X sky130_fd_sc_hd__mux2_1
XFILLER_3_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10305_ VGND VPWR VPWR VGND _10305_/X hold374/A _11098_/S hold606/A sky130_fd_sc_hd__mux2_1
X_11285_ VGND VPWR VPWR VGND _11286_/B _14811_/Q _11299_/S _14379_/Q sky130_fd_sc_hd__mux2_1
X_10236_ VGND VPWR VGND VPWR _10236_/X _11235_/A1 _10232_/X _10235_/X _11235_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_80_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10167_ VGND VPWR VPWR VGND _10167_/X _10166_/X _10467_/S _10165_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14975_ hold412/A _14975_/CLK _14975_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10098_ VPWR VGND VPWR VGND _10097_/X _10608_/A1 _10096_/X _10098_/Y sky130_fd_sc_hd__a21oi_1
X_13278__395 VPWR VGND VPWR VGND _14553_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_12808_ VGND VPWR VPWR VGND _12809_/B _07962_/Y _12820_/B _07959_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1093 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12739_ VGND VPWR VGND VPWR _12739_/X _12738_/X _12737_/X _12735_/S _12739_/C1 sky130_fd_sc_hd__a211o_1
X_15527_ hold300/A _15527_/CLK _15527_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15458_ _15458_/Q clkload16/A _15458_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14409_ _14409_/Q clkload39/A _14409_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_15389_ hold687/A _15389_/CLK _15389_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold526 hold526/X hold526/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 hold515/X hold515/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 hold504/X hold504/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ VPWR VGND VPWR VGND _09949_/Y hold1322/X _09956_/S _14128_/D _09937_/Y sky130_fd_sc_hd__a22o_1
Xhold559 hold559/X hold559/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 hold537/X hold537/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 hold548/X hold548/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08901_ VGND VPWR VGND VPWR _15142_/D hold1339/X _08902_/B _08900_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
X_09881_ VPWR VGND VPWR VGND _09877_/X hold226/X _09880_/Y _09882_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08832_ VGND VPWR VPWR VGND _15181_/D fanout38/X _08844_/S hold726/X sky130_fd_sc_hd__mux2_1
XFILLER_44_1048 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_39_920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1204 hold1204/X _14465_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 hold1215/X _14265_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _09894_/S _14146_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08763_ VGND VPWR VPWR VGND _15243_/D fanout32/X _08779_/S hold231/X sky130_fd_sc_hd__mux2_1
Xhold1248 hold1248/X _14625_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 hold1226/X _14891_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07714_ VPWR VGND _07714_/A _07714_/X _07826_/D VPWR VGND sky130_fd_sc_hd__and2_2
Xhold1259 hold1259/X _14334_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13519__636 VPWR VGND VPWR VGND _14794_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
XFILLER_2_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08694_ VGND VPWR VGND VPWR _08694_/X _08700_/A2 _08700_/B1 hold978/X _08693_/X sky130_fd_sc_hd__a211o_1
X_07645_ VPWR VGND VPWR VGND _15132_/Q clone19/X _15359_/Q clone13/X _07645_/X sky130_fd_sc_hd__a22o_2
X_07576_ VGND VPWR VGND VPWR _07575_/Y _07523_/Y _07487_/B _08591_/B _09007_/B _15547_/Q
+ sky130_fd_sc_hd__a32oi_4
X_14117__1234 VPWR VGND VPWR VGND _15536_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_09315_ VGND VPWR VPWR VGND _14729_/D hold911/X _09342_/S clone133/X sky130_fd_sc_hd__mux2_1
XFILLER_55_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09246_ VGND VPWR VPWR VGND _14797_/D clone45/X _09269_/S hold732/X sky130_fd_sc_hd__mux2_1
XFILLER_22_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_31_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09177_ VGND VPWR VPWR VGND _14914_/D hold387/X _09194_/S fanout44/X sky130_fd_sc_hd__mux2_1
XFILLER_31_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08128_ VGND VPWR VGND VPWR _08127_/X fanout7/A _08128_/A _08128_/B sky130_fd_sc_hd__or3b_4
X_13071__188 VPWR VGND VPWR VGND _14314_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_08059_ VGND VPWR _08059_/B _08060_/B _15555_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_11070_ VGND VPWR VGND VPWR _11070_/X _11181_/A1 _11065_/X _11069_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
X_10021_ VPWR VGND VGND VPWR _10021_/A _10021_/B _10022_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_40_1424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14760_ hold299/A _14760_/CLK _14760_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11972_ VPWR VGND VGND VPWR _11953_/X _11970_/X _07913_/Y _11971_/X _11972_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14001__1118 VPWR VGND VPWR VGND _15373_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_14691_ hold754/A _14691_/CLK _14691_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10923_ VGND VPWR VPWR VGND _10923_/X hold610/A _11240_/S hold288/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_73_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10854_ VGND VPWR VGND VPWR _10854_/X _10851_/A _10850_/X _10853_/X _11096_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_73_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15312_ hold886/A _15312_/CLK _15312_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10785_ VPWR VGND VGND VPWR _10766_/Y _10784_/X _12269_/B _14397_/Q _14397_/D _11341_/A
+ sky130_fd_sc_hd__o221a_1
X_12524_ VPWR VGND VGND VPWR _12524_/X hold358/A _12736_/B sky130_fd_sc_hd__or2_1
X_13312__429 VPWR VGND VPWR VGND _14587_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_12_374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15243_ hold231/A _15243_/CLK _15243_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12455_ VPWR VGND VGND VPWR _12436_/Y _12454_/X _12677_/A2 _15468_/Q _15468_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_11406_ VGND VPWR _11406_/X _11410_/A _14856_/Q _11406_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_13930__1047 VPWR VGND VPWR VGND _15302_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_12386_ VPWR VGND VGND VPWR _12386_/X _12721_/S _12386_/B sky130_fd_sc_hd__or2_1
X_15174_ hold367/A _15174_/CLK _15174_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12906__23 VPWR VGND VPWR VGND _14148_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_11337_ VPWR VGND VGND VPWR _11336_/Y _11421_/C _11316_/Y _14831_/Q _14831_/D _11337_/C1
+ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13663__780 VPWR VGND VPWR VGND _15003_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_11268_ VPWR VGND VGND VPWR _11269_/B _15431_/Q _11541_/B sky130_fd_sc_hd__or2_1
X_13206__323 VPWR VGND VPWR VGND _14481_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_11199_ VGND VPWR VPWR VGND _11199_/X _11196_/X _11213_/S _11195_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10219_ VGND VPWR VGND VPWR _10219_/X _11237_/A1 _10214_/X _10218_/X _12869_/A1 sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_36_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14958_ hold961/A _14958_/CLK _14958_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14889_ _14889_/Q _14889_/CLK _14889_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_915 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_35_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07430_ VPWR VGND VGND VPWR _15465_/Q _07512_/A _07511_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_56_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07361_ VPWR VGND VPWR VGND _08290_/B _07229_/A _08278_/A _08275_/A _08290_/A sky130_fd_sc_hd__a22o_1
X_09100_ VGND VPWR VPWR VGND _14995_/D hold263/X _09124_/S fanout77/X sky130_fd_sc_hd__mux2_1
X_07292_ VPWR VGND VGND VPWR _07293_/B _15468_/Q _07292_/B sky130_fd_sc_hd__or2_1
X_09031_ VGND VPWR VPWR VGND _15059_/D hold655/X _09055_/S fanout77/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold301 hold301/X hold301/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 hold323/X hold323/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 hold334/X hold334/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 hold312/X hold312/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 hold356/X hold356/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 hold378/X hold378/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 hold367/X hold367/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 hold345/X hold345/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout825 VPWR VGND _09024_/A _09977_/A VPWR VGND sky130_fd_sc_hd__buf_2
X_09933_ VPWR VGND VGND VPWR hold539/X _09931_/Y _09932_/Y _14133_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout814 VPWR VGND _12159_/C1 fanout829/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout803 VGND VPWR _11296_/A _11290_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold389 hold389/X hold389/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout836 VPWR VGND _09976_/B fanout844/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_63_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout847 VGND VPWR _07422_/X _08263_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09864_ VGND VPWR VPWR VGND _14158_/D hold439/X _09864_/S _09864_/A0 sky130_fd_sc_hd__mux2_1
Xhold1012 _15121_/D _08951_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1023 hold1023/X _14349_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ VPWR VGND VGND VPWR _09095_/B _09556_/C _09240_/A _09311_/B sky130_fd_sc_hd__nand3b_1
Xfanout869 VPWR VGND _07519_/B _07511_/B VPWR VGND sky130_fd_sc_hd__buf_2
Xhold1001 hold1001/X _14489_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1056 hold1056/X _15108_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1045 hold1045/X _14501_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 hold1034/X _15294_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ VGND VPWR VPWR VGND _14254_/D _09864_/A0 _09795_/S hold492/X sky130_fd_sc_hd__mux2_1
XFILLER_6_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1067 hold1067/X _14876_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 hold1089/X _14450_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1078 hold1078/X _15012_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ VPWR VGND VPWR VGND _08746_/Y _08776_/S sky130_fd_sc_hd__inv_2
X_08677_ VGND VPWR VGND VPWR _15289_/D hold1100/X _08686_/A2 _08676_/X _12085_/C1
+ sky130_fd_sc_hd__o211a_1
X_07628_ _07629_/C _07624_/X _07625_/Y _07627_/X _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_26_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07559_ VPWR VGND VPWR VGND _07560_/B _07560_/C _11284_/A _07559_/A _07560_/D sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_64_Right_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10570_ VGND VPWR VPWR VGND _10570_/X _10567_/X _10732_/S _10566_/X sky130_fd_sc_hd__mux2_1
X_09229_ VGND VPWR VPWR VGND _14864_/D hold927/X _09229_/S _09229_/A0 sky130_fd_sc_hd__mux2_1
X_13647__764 VPWR VGND VPWR VGND _14987_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_12240_ VGND VPWR VPWR VGND _12240_/X hold479/A _12318_/S hold256/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12171_ VGND VPWR VPWR VGND _12171_/X hold694/A _12171_/S hold242/A sky130_fd_sc_hd__mux2_1
Xhold890 hold890/X hold890/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11122_ VGND VPWR VPWR VGND _11122_/X hold456/A _11142_/S hold326/A sky130_fd_sc_hd__mux2_1
X_11053_ VGND VPWR VPWR VGND _11057_/B hold641/A _11165_/S hold283/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10004_ VPWR VGND VPWR VGND _10003_/C _15616_/Q hold1309/X _10005_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14812_ _14812_/Q clkload20/A _14812_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_64_528 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11955_ VGND VPWR VPWR VGND _11958_/B hold929/A _11964_/S hold572/A sky130_fd_sc_hd__mux2_1
X_14743_ hold659/A _14743_/CLK _14743_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14674_ hold435/A _14674_/CLK _14674_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10906_ VGND VPWR VPWR VGND _10906_/X _14273_/Q _10919_/S _14305_/Q sky130_fd_sc_hd__mux2_1
X_11886_ VGND VPWR VPWR VGND _11886_/X _11883_/X _12164_/A _11882_/X sky130_fd_sc_hd__mux2_1
X_10837_ VGND VPWR VGND VPWR _10837_/X _10834_/X _10836_/X _11086_/C1 _11218_/A1 sky130_fd_sc_hd__a211o_1
X_10768_ VGND VPWR VPWR VGND _10768_/X hold869/A _11091_/S hold742/A sky130_fd_sc_hd__mux2_1
XFILLER_41_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12507_ VGND VPWR VPWR VGND _12507_/X _12504_/X _12536_/S _12503_/X sky130_fd_sc_hd__mux2_1
X_10699_ VGND VPWR VPWR VGND _10703_/B hold705/A _10700_/S hold420/A sky130_fd_sc_hd__mux2_1
X_12438_ VGND VPWR VPWR VGND _12438_/X hold866/A _12661_/S hold454/A sky130_fd_sc_hd__mux2_1
X_15226_ _15226_/Q _15226_/CLK _15226_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15157_ _15157_/Q _15157_/CLK _15157_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12369_ VGND VPWR VPWR VGND _12373_/B _15184_/Q _12370_/S hold707/A sky130_fd_sc_hd__mux2_1
X_15088_ _15088_/Q clkload36/A _15088_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_79_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14214__932 _14214_/D _14214__932/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_14116__1233 VPWR VGND VPWR VGND _15535_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_13440__557 VPWR VGND VPWR VGND _14715_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_80_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08600_ VPWR VGND VGND VPWR _08605_/A _08998_/B _08600_/Y sky130_fd_sc_hd__nor2_1
X_09580_ VGND VPWR VPWR VGND _14485_/D hold1015/X _09590_/S fanout9/X sky130_fd_sc_hd__mux2_1
X_08531_ VPWR VGND _15321_/D _08531_/B _11398_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_36_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13293__410 VPWR VGND VPWR VGND _14568_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_08462_ VPWR VGND VGND VPWR _08462_/X _15345_/Q _08482_/B sky130_fd_sc_hd__or2_1
X_07413_ VPWR VGND VPWR VGND _07413_/Y _07412_/X _07333_/Y _07326_/Y _07329_/X sky130_fd_sc_hd__a211oi_1
XFILLER_1_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13334__451 VPWR VGND VPWR VGND _14609_/CLK clkload52/A sky130_fd_sc_hd__inv_2
X_08393_ VGND VPWR VPWR VGND _15384_/D fanout38/X _08393_/S hold599/X sky130_fd_sc_hd__mux2_1
X_07344_ _07389_/A _07876_/A _07820_/A _07859_/A _07899_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_32_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07275_ VPWR VGND VGND VPWR _07981_/B _07981_/A _07971_/A _07916_/A sky130_fd_sc_hd__nor3_1
XFILLER_17_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09014_ VGND VPWR VGND VPWR _09014_/X _09873_/A _09016_/B1 _15098_/Q _09013_/Y sky130_fd_sc_hd__a211o_1
XFILLER_30_1412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold153 hold153/X hold153/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14000__1117 VPWR VGND VPWR VGND _15372_/CLK clkload55/A sky130_fd_sc_hd__inv_2
Xhold175 hold175/X hold175/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/X hold186/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/X hold164/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ VGND VPWR VPWR VGND _09916_/A _09917_/B _09916_/B sky130_fd_sc_hd__xor2_1
X_12897__14 VPWR VGND VPWR VGND _14139_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
Xfanout611 VPWR VGND _08231_/S _08251_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout622 VPWR VGND _09864_/S _09834_/Y VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout633 VPWR VGND _09687_/S _09690_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xhold197 hold197/X hold197/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 VPWR VGND _08779_/S _08772_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout655 VPWR VGND _09467_/S _09482_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout644 VPWR VGND _09555_/S _09553_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout666 VPWR VGND _09229_/S _09198_/X VPWR VGND sky130_fd_sc_hd__buf_4
X_09847_ VGND VPWR VPWR VGND _14175_/D hold767/X _09861_/S fanout46/X sky130_fd_sc_hd__mux2_1
Xfanout677 VGND VPWR _09095_/X _09125_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout699 VGND VPWR _12877_/S _12860_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout688 VGND VPWR _08304_/X _08330_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09778_ VGND VPWR VPWR VGND _14271_/D fanout46/X _09795_/S hold970/X sky130_fd_sc_hd__mux2_1
XFILLER_37_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08729_ VGND VPWR VGND VPWR _15269_/D hold1020/X _08731_/A2 _08728_/X _11294_/A sky130_fd_sc_hd__o211a_1
XFILLER_2_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11740_ VGND VPWR VGND VPWR _11740_/X _11739_/X _11738_/X _12396_/S _12720_/C1 sky130_fd_sc_hd__a211o_1
X_11671_ VGND VPWR VGND VPWR _11671_/X _11668_/X _11670_/X _11894_/S _12189_/C1 sky130_fd_sc_hd__a211o_1
X_13077__194 VPWR VGND VPWR VGND _14320_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_14390_ _14390_/Q clkload11/A _14390_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10622_ VGND VPWR VGND VPWR _10622_/X _10621_/X _10620_/X _10634_/A1 _10622_/C1 sky130_fd_sc_hd__a211o_1
X_10553_ VGND VPWR VPWR VGND _10553_/X hold902/A _10553_/S hold352/A sky130_fd_sc_hd__mux2_1
X_13881__998 VPWR VGND VPWR VGND _15253_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_10484_ VPWR VGND VGND VPWR _10484_/X hold391/A _10484_/B sky130_fd_sc_hd__or2_1
X_15011_ hold995/A _15011_/CLK _15011_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12223_ VGND VPWR VPWR VGND _12223_/X hold633/A _12227_/S hold266/A sky130_fd_sc_hd__mux2_1
X_12154_ VGND VPWR VGND VPWR _12154_/X hold936/A _12229_/A2 _12147_/S _12153_/X sky130_fd_sc_hd__o211a_1
X_11105_ VPWR VGND VPWR VGND _11102_/X _11112_/A _11104_/X _11105_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_620 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12085_ VPWR VGND VGND VPWR _12066_/Y _12084_/X _12380_/B _15458_/Q _15458_/D _12085_/C1
+ sky130_fd_sc_hd__o221a_1
XFILLER_77_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11036_ VGND VPWR VGND VPWR _11036_/X _15024_/Q _11252_/A2 _11035_/X _11250_/S sky130_fd_sc_hd__o211a_1
XFILLER_65_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13775__892 VPWR VGND VPWR VGND _15147_/CLK clkload32/A sky130_fd_sc_hd__inv_2
XFILLER_40_1073 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14726_ _14726_/Q _14726_/CLK _14726_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11938_ VGND VPWR VPWR VGND _11938_/X hold554/A _11950_/B hold607/A sky130_fd_sc_hd__mux2_1
X_13318__435 VPWR VGND VPWR VGND _14593_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XFILLER_53_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11869_ VGND VPWR VGND VPWR _11869_/X hold884/A _12192_/A2 _11958_/A _11868_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14657_ hold450/A _14657_/CLK _14657_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_60_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14588_ hold237/A _14588_/CLK _14588_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12991__108 VPWR VGND VPWR VGND _14234_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_14_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15209_ _15209_/Q _15209_/CLK _15209_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12981__98 VPWR VGND VPWR VGND _14224_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_09701_ VGND VPWR VPWR VGND _14342_/D _09710_/S clone47/X hold1271/X sky130_fd_sc_hd__mux2_4
X_07962_ VPWR VGND VGND VPWR _07962_/A _07962_/B _07962_/Y sky130_fd_sc_hd__nor2_1
X_07893_ VGND VPWR VPWR VGND _07893_/X _07558_/A _08902_/A _07567_/B _07892_/Y sky130_fd_sc_hd__o31a_4
X_09632_ VGND VPWR VPWR VGND _14438_/D _09637_/S hold1199/X clone111/X sky130_fd_sc_hd__mux2_4
X_09563_ VGND VPWR VPWR VGND _14502_/D _09584_/S hold1177/X fanout74/X sky130_fd_sc_hd__mux2_4
X_08514_ VPWR VGND _15329_/D _08514_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
X_09494_ VGND VPWR VPWR VGND _14565_/D fanout70/X _09517_/S hold695/X sky130_fd_sc_hd__mux2_1
X_08445_ VGND VPWR VGND VPWR _15354_/D hold1398/X _08448_/B _08444_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_12_918 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08376_ VPWR VGND VPWR VGND _15577_/Q _09198_/B _09164_/A _09694_/A sky130_fd_sc_hd__or3_4
X_07327_ VPWR VGND _07327_/X _07328_/B _11535_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_13111__228 VPWR VGND VPWR VGND _14354_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_07258_ VPWR VGND _07271_/B _07258_/B _15458_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07189_ VPWR VGND VGND VPWR _07190_/B _15456_/Q _07189_/B sky130_fd_sc_hd__or2_1
XFILLER_2_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout441 VGND VPWR _07851_/Y _11023_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13759__876 VPWR VGND VPWR VGND _15131_/CLK clkload23/A sky130_fd_sc_hd__inv_2
Xfanout430 VGND VPWR _10505_/A1 _10667_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout452 VGND VPWR _12869_/A1 _11218_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout474 VPWR VGND VGND VPWR _07569_/X _12080_/A2 sky130_fd_sc_hd__buf_12
XFILLER_58_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout463 VGND VPWR _12118_/A2 _12040_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout496 VGND VPWR fanout497/X _11965_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout485 VGND VPWR _12005_/S _12112_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_62_807 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12841_ VGND VPWR VGND VPWR _15569_/D _07222_/A _11458_/S _11480_/S _12840_/Y sky130_fd_sc_hd__o211a_1
XFILLER_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13005__122 VPWR VGND VPWR VGND _14248_/CLK clkload41/A sky130_fd_sc_hd__inv_2
XFILLER_73_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12772_ VPWR VGND VGND VPWR _12772_/A _12788_/S _12772_/Y sky130_fd_sc_hd__nor2_1
X_15560_ _15560_/Q clkload44/A _15560_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15491_ _15491_/Q _15491_/CLK _15491_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11723_ VPWR VGND VPWR VGND _11722_/X _12415_/C1 _11721_/X _11723_/Y sky130_fd_sc_hd__a21oi_1
X_14511_ hold167/A _14511_/CLK _14511_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14115__1232 VPWR VGND VPWR VGND _15534_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_11654_ VPWR VGND VGND VPWR _11654_/X _11948_/S _11654_/B sky130_fd_sc_hd__or2_1
XFILLER_42_575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14442_ _14442_/Q _14442_/CLK _14442_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout70 VGND VPWR fanout71/X fanout70/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout92 VPWR VGND fanout92/X fanout93/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout81 VPWR VGND VGND VPWR clone49/A fanout81/X sky130_fd_sc_hd__buf_8
X_10605_ VPWR VGND VGND VPWR _10605_/X _10613_/A _10605_/B sky130_fd_sc_hd__or2_1
X_14373_ hold783/A _14373_/CLK _14373_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11585_ VPWR VGND VGND VPWR _12103_/A _11585_/B _11585_/Y sky130_fd_sc_hd__nor2_1
X_10536_ VGND VPWR VPWR VGND _10536_/X _14455_/Q _10700_/S hold659/A sky130_fd_sc_hd__mux2_1
XFILLER_10_483 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10467_ VGND VPWR VPWR VGND _10467_/X _10464_/X _10467_/S _10463_/X sky130_fd_sc_hd__mux2_1
X_13703__820 VPWR VGND VPWR VGND _15043_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_12206_ VGND VPWR VPWR VGND _12206_/X hold544/A _12228_/B hold408/A sky130_fd_sc_hd__mux2_1
X_10398_ VGND VPWR VPWR VGND _10398_/X hold861/A _10696_/S hold710/A sky130_fd_sc_hd__mux2_1
X_12137_ VGND VPWR VPWR VGND _12137_/X _12134_/X _12147_/S _12133_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12068_ VGND VPWR VPWR VGND _12068_/X hold857/A _12219_/S hold634/A sky130_fd_sc_hd__mux2_1
X_11019_ VGND VPWR VPWR VGND _11019_/X hold587/A _11165_/S hold441/A sky130_fd_sc_hd__mux2_1
X_13552__669 VPWR VGND VPWR VGND _14883_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_14709_ hold572/A _14709_/CLK _14709_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08230_ VPWR VGND VPWR VGND _08220_/X _08230_/X _08230_/A _08230_/B sky130_fd_sc_hd__or3b_2
X_08161_ VGND VPWR _07372_/C _08181_/A _08162_/B _07372_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_07112_ VPWR VGND VPWR VGND _07827_/A _07703_/A sky130_fd_sc_hd__inv_2
X_08092_ VGND VPWR VPWR VGND _15524_/D fanout13/X _08300_/S hold216/X sky130_fd_sc_hd__mux2_1
Xclkload51 VGND VPWR VPWR VGND clkload51/A clkload51/Y sky130_fd_sc_hd__clkinv_2
Xclkload40 VGND VPWR VPWR VGND clkload40/A clkload40/Y sky130_fd_sc_hd__clkinvlp_4
X_13446__563 VPWR VGND VPWR VGND _14721_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_08994_ VGND VPWR VGND VPWR _15106_/D hold1031/X _09015_/A2 _08993_/X _09000_/C1
+ sky130_fd_sc_hd__o211a_1
X_07945_ VPWR VGND VGND VPWR _07945_/A _10075_/A _07945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_1322 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09615_ VGND VPWR VPWR VGND _14453_/D fanout8/X _09625_/S hold596/X sky130_fd_sc_hd__mux2_1
X_07876_ VGND VPWR _07876_/B _12826_/B _07876_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_3_1195 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09546_ VGND VPWR VPWR VGND _14516_/D fanout5/X _09555_/S hold158/X sky130_fd_sc_hd__mux2_1
X_09477_ VGND VPWR VPWR VGND _14579_/D _09859_/A0 _09485_/S hold178/X sky130_fd_sc_hd__mux2_1
X_08428_ VPWR VGND VGND VPWR _08428_/X _08428_/A _08484_/B sky130_fd_sc_hd__or2_1
XFILLER_71_1331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 VPWR VGND VPWR VGND clkload1/Y clkload1/A sky130_fd_sc_hd__inv_6
X_08359_ VGND VPWR VPWR VGND _15414_/D hold380/X _08366_/S fanout33/X sky130_fd_sc_hd__mux2_1
X_11370_ VGND VPWR VPWR VGND _14843_/D _11369_/X _11382_/S hold1404/X sky130_fd_sc_hd__mux2_1
X_10321_ VGND VPWR VPWR VGND _10321_/X hold962/A _11261_/B hold397/A sky130_fd_sc_hd__mux2_1
XFILLER_4_903 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10252_ VGND VPWR VGND VPWR _10252_/X _10251_/X _10250_/X _11235_/A1 _10918_/C1 sky130_fd_sc_hd__a211o_1
X_10183_ VGND VPWR VPWR VGND _10187_/B hold809/A _10479_/S hold188/A sky130_fd_sc_hd__mux2_1
X_14991_ hold301/A _14991_/CLK _14991_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout260 VPWR VGND _12583_/S _12694_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout282 VPWR VGND fanout282/X _07894_/X VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_47_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout271 VGND VPWR _10629_/A2 _10633_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout293 VGND VPWR _10520_/S _10627_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_35_807 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12824_ VPWR VGND VGND VPWR _12822_/Y _12823_/X _15563_/Q _10056_/A _15563_/D _07544_/B
+ sky130_fd_sc_hd__o221a_1
X_15612_ _15612_/Q clkload27/A _15612_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12755_ VPWR VGND VGND VPWR _08246_/Y _10079_/X _08240_/B _12789_/A _12755_/X _10060_/A
+ sky130_fd_sc_hd__o221a_1
X_15543_ hold325/A _15543_/CLK _15543_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_30_512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11706_ VPWR VGND VGND VPWR _11706_/X hold275/A _12716_/S sky130_fd_sc_hd__or2_1
X_12686_ VGND VPWR VPWR VGND _12690_/B hold489/A _12689_/S hold377/A sky130_fd_sc_hd__mux2_1
X_15474_ _15474_/Q clkload40/A _15474_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13389__506 VPWR VGND VPWR VGND _14664_/CLK clkload41/A sky130_fd_sc_hd__inv_2
XFILLER_30_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11637_ VGND VPWR VGND VPWR _11637_/X _15000_/Q _12040_/A2 _11625_/S _11636_/X sky130_fd_sc_hd__o211a_1
X_14425_ hold800/A _14425_/CLK _14425_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13133__250 VPWR VGND VPWR VGND _14376_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_11568_ VGND VPWR VPWR VGND _11572_/B hold876/A _12094_/S hold692/A sky130_fd_sc_hd__mux2_1
X_14356_ hold981/A _14356_/CLK _14356_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold708 hold708/X hold708/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ VGND VPWR VGND VPWR _10519_/X _10516_/X _10518_/X _10523_/A1 _10630_/C1 sky130_fd_sc_hd__a211o_1
Xhold719 hold719/X hold719/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11499_ VGND VPWR VPWR VGND _11499_/X _15085_/Q _11535_/C _15083_/Q sky130_fd_sc_hd__mux2_1
X_14287_ hold255/A _14287_/CLK _14287_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12951__68 VPWR VGND VPWR VGND _14194_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
Xhold1408 hold1408/X _14931_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07730_ VGND VPWR VPWR VGND _15558_/Q _07798_/A _07730_/B sky130_fd_sc_hd__xor2_1
Xhold1419 _07082_/A _15567_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07661_ VPWR VGND VPWR VGND _15131_/Q _07873_/B1 _15358_/Q _07558_/B _07661_/X sky130_fd_sc_hd__a22o_2
X_12997__114 VPWR VGND VPWR VGND _14240_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_07592_ VGND VPWR VGND VPWR _15355_/Q _08495_/A2 _07873_/B1 _07592_/Y _15144_/Q sky130_fd_sc_hd__a22oi_4
XFILLER_53_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09400_ VGND VPWR VPWR VGND _14649_/D hold667/X _09414_/S fanout23/X sky130_fd_sc_hd__mux2_1
XFILLER_19_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09331_ VGND VPWR VPWR VGND _14713_/D hold724/X _09345_/S fanout26/X sky130_fd_sc_hd__mux2_1
XFILLER_34_884 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09262_ VGND VPWR VPWR VGND _14781_/D fanout19/X _09268_/S hold574/X sky130_fd_sc_hd__mux2_1
XFILLER_21_534 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08213_ VGND VPWR VPWR VGND _15518_/D _09550_/A1 _08300_/S hold314/X sky130_fd_sc_hd__mux2_1
X_09193_ VGND VPWR VPWR VGND _14898_/D hold578/X _09194_/S _09689_/A0 sky130_fd_sc_hd__mux2_1
X_08144_ VPWR VGND VGND VPWR _15551_/Q _08155_/A _08145_/B sky130_fd_sc_hd__nor2_1
XFILLER_66_1411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08075_ VPWR VGND VGND VPWR _07574_/A _08074_/X _07996_/X _08075_/X sky130_fd_sc_hd__o21a_1
X_13680__797 VPWR VGND VPWR VGND _15020_/CLK clkload45/A sky130_fd_sc_hd__inv_2
XFILLER_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08977_ VPWR VGND VGND VPWR _08983_/A _08977_/B _08977_/Y sky130_fd_sc_hd__nor2_1
X_14114__1231 VPWR VGND VPWR VGND _15533_/CLK clkload53/A sky130_fd_sc_hd__inv_2
XFILLER_29_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_1213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_9_1382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07928_ _07933_/B _07924_/X _07925_/Y _07927_/X _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07859_ VPWR VGND VGND VPWR _07859_/A _07859_/B _07859_/Y sky130_fd_sc_hd__nor2_1
X_10870_ VGND VPWR VPWR VGND _10870_/X _10869_/X _11110_/A _10868_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13574__691 VPWR VGND VPWR VGND _14905_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
XFILLER_16_328 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09529_ VGND VPWR VPWR VGND _14533_/D fanout68/X _09549_/S hold157/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12540_ VGND VPWR VPWR VGND _12540_/X _14213_/Q _12652_/S hold285/A sky130_fd_sc_hd__mux2_1
XFILLER_40_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12471_ VPWR VGND VPWR VGND _12470_/X _12722_/A1 _12469_/X _12471_/Y sky130_fd_sc_hd__a21oi_1
X_13117__234 VPWR VGND VPWR VGND _14360_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_11422_ VGND VPWR VGND VPWR _11422_/X _14926_/Q _11303_/A _11431_/A2 sky130_fd_sc_hd__a21bo_1
X_15190_ hold691/A _15190_/CLK _15190_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14210_ _14210_/Q _14210_/CLK _14210_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14141_ hold819/A _14141_/CLK _14141_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11353_ VGND VPWR VPWR VGND _11353_/X _14931_/Q _11355_/S hold1187/X sky130_fd_sc_hd__mux2_1
XFILLER_10_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11284_ VGND VPWR VGND VPWR _11302_/B _11299_/S _11284_/A _11284_/B sky130_fd_sc_hd__or3b_4
XFILLER_10_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10304_ VPWR VGND VGND VPWR _10285_/Y _10303_/X _10192_/B _14384_/Q _14384_/D _12159_/C1
+ sky130_fd_sc_hd__o221a_1
X_10235_ VPWR VGND VGND VPWR _10235_/X _10911_/S _10235_/B sky130_fd_sc_hd__or2_1
X_10166_ VGND VPWR VPWR VGND _10166_/X hold681/A _10169_/B hold297/A sky130_fd_sc_hd__mux2_1
XFILLER_67_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14974_ hold524/A _14974_/CLK _14974_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10097_ VGND VPWR VPWR VGND _10097_/X _10094_/X _10613_/A _10093_/X sky130_fd_sc_hd__mux2_1
X_13815__932 VPWR VGND VPWR VGND _15187_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_12807_ VGND VPWR VPWR VGND _15559_/D _12806_/Y _12805_/Y _12807_/A1 _12807_/B1 _15559_/Q
+ sky130_fd_sc_hd__a32o_1
X_10999_ VGND VPWR VGND VPWR _10999_/X _15505_/Q _11003_/A2 _10998_/X _10985_/S sky130_fd_sc_hd__o211a_1
XFILLER_42_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12738_ VGND VPWR VPWR VGND _12738_/X _14893_/Q _12747_/S _15429_/Q sky130_fd_sc_hd__mux2_1
X_15526_ hold238/A _15526_/CLK _15526_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15457_ _15457_/Q clkload13/A _15457_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12669_ VGND VPWR VGND VPWR _12669_/X hold959/A _12669_/A2 _12735_/S _12668_/X sky130_fd_sc_hd__o211a_1
XFILLER_15_1354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14408_ _14408_/Q clkload40/A _14408_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_15388_ hold610/A _15388_/CLK _15388_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold505 hold505/X hold505/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 hold527/X hold527/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14339_ hold482/A _14339_/CLK _14339_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold516 hold516/X hold516/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 hold549/X hold549/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 hold538/X hold538/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09880_ VPWR VGND VGND VPWR _09885_/C _09880_/B _09880_/Y sky130_fd_sc_hd__nor2_1
X_08900_ VPWR VGND VGND VPWR _08900_/X _15142_/Q _08924_/B sky130_fd_sc_hd__or2_1
XFILLER_48_1141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_48_1196 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08831_ VGND VPWR VPWR VGND _15182_/D fanout41/X _08844_/S hold853/X sky130_fd_sc_hd__mux2_1
Xhold1216 hold1216/X _15324_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1205 hold1205/X _15359_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 _11273_/A _15436_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 hold1249/X _15153_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ VGND VPWR VPWR VGND _15244_/D fanout36/X _08772_/S hold258/X sky130_fd_sc_hd__mux2_1
Xhold1227 hold1227/X _14344_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13558__675 VPWR VGND VPWR VGND _14889_/CLK clkload47/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_69_Left_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_66_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_1396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07713_ VPWR VGND VGND VPWR _15563_/Q _07803_/B _07713_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08693_ VGND VPWR VGND VPWR _08693_/X _14394_/Q _08640_/B _08711_/B1 _08629_/X sky130_fd_sc_hd__o211a_1
XFILLER_39_998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07644_ VGND VPWR VPWR VGND _15541_/D fanout77/X _08231_/S hold164/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07575_ VGND VPWR _07575_/A2 _07486_/A _07575_/Y _07486_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_15_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09314_ _14730_/D fanout92/X fanout88/X _09327_/S _09313_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09245_ VGND VPWR VPWR VGND _14798_/D fanout84/X _09272_/S hold489/X sky130_fd_sc_hd__mux2_1
X_09176_ VGND VPWR VPWR VGND _09194_/S hold1081/X fanout50/X _14915_/D sky130_fd_sc_hd__mux2_2
X_08127_ VGND VPWR VPWR VGND _08127_/X _07996_/X _08114_/Y _08147_/A _12776_/A sky130_fd_sc_hd__o2bb2a_1
X_08058_ VPWR VGND VGND VPWR _08147_/A _08058_/B _08070_/B sky130_fd_sc_hd__nor2_1
X_14190__908 _14190_/D _14190__908/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_10020_ VPWR VGND _10024_/C _10021_/B _15624_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_11971_ VPWR VGND _11971_/X _11945_/X _11941_/X _12111_/C1 _12029_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_57_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_5_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10922_ VGND VPWR VGND VPWR _10922_/X _10930_/C1 _10921_/X _10918_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
X_14690_ hold991/A _14690_/CLK _14690_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10853_ VPWR VGND VGND VPWR _10853_/X _11112_/A _10853_/B sky130_fd_sc_hd__or2_1
X_10784_ VPWR VGND VPWR VGND _10783_/X _07691_/X _12602_/B1 _10784_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15311_ _15311_/Q _15311_/CLK _15311_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12523_ VGND VPWR VPWR VGND _12523_/X hold775/A _12736_/B hold527/A sky130_fd_sc_hd__mux2_1
X_15242_ hold273/A _15242_/CLK _15242_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13351__468 VPWR VGND VPWR VGND _14626_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_12454_ VPWR VGND VPWR VGND _12453_/X _12658_/A _12713_/B1 _12454_/X sky130_fd_sc_hd__a21o_1
X_11405_ VGND VPWR VGND VPWR _14855_/D _14855_/Q _11408_/A _11404_/Y _08541_/A sky130_fd_sc_hd__o211a_1
X_15173_ hold794/A _15173_/CLK _15173_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12385_ VGND VPWR VPWR VGND _12385_/X _14561_/Q _12408_/S _14593_/Q sky130_fd_sc_hd__mux2_1
X_11336_ VPWR VGND VGND VPWR _11338_/B _11336_/B _11336_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_1450 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11267_ VPWR VGND VGND VPWR _11541_/B _15430_/Q _14800_/Q sky130_fd_sc_hd__or2_1
XFILLER_45_1325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11198_ VGND VPWR VGND VPWR _11198_/X _11215_/C1 _11194_/X _11197_/X _11217_/C1 sky130_fd_sc_hd__o211a_1
X_12921__38 VPWR VGND VPWR VGND _14164_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_13245__362 VPWR VGND VPWR VGND _14520_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_10218_ VGND VPWR VGND VPWR _10218_/X _10217_/X _10216_/X _10995_/S _11235_/C1 sky130_fd_sc_hd__a211o_1
X_10149_ VGND VPWR VGND VPWR _10149_/X _10146_/X _10148_/X _10523_/A1 _10630_/C1 sky130_fd_sc_hd__a211o_1
X_14957_ hold831/A _14957_/CLK _14957_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14888_ hold935/A _14888_/CLK _14888_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_50_448 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07360_ VPWR VGND VGND VPWR _08258_/B _07360_/A _07360_/B sky130_fd_sc_hd__or2_1
X_15509_ hold824/A _15509_/CLK _15509_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14113__1230 VPWR VGND VPWR VGND _15532_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_07291_ VPWR VGND _07291_/X _07292_/B _15468_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_09030_ VGND VPWR VPWR VGND _15060_/D hold624/X _09055_/S fanout80/X sky130_fd_sc_hd__mux2_1
Xhold302 hold302/X hold302/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 hold324/X hold324/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 hold313/X hold313/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/X hold335/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ VPWR VGND VPWR VGND _09931_/Y hold539/X _09917_/A _09932_/Y sky130_fd_sc_hd__a21oi_1
Xhold357 hold357/X hold357/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 hold368/X hold368/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 hold346/X hold346/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 hold379/X hold379/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout804 VPWR VGND _11296_/A fanout829/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout815 VPWR VGND _11937_/C1 _12233_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout837 VPWR VGND _08955_/A _08943_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout826 VPWR VGND _09977_/A _08571_/B VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout848 VGND VPWR _07422_/X _10074_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09863_ VGND VPWR VPWR VGND _14159_/D hold731/X _09864_/S _09863_/A0 sky130_fd_sc_hd__mux2_1
Xhold1013 hold1013/X _14545_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout859 VPWR VGND _10059_/A _07137_/X VPWR VGND sky130_fd_sc_hd__buf_6
X_08814_ VGND VPWR VPWR VGND _15195_/D fanout97/X _08814_/S hold224/X sky130_fd_sc_hd__mux2_1
X_09794_ VGND VPWR VPWR VGND _14255_/D _09829_/A1 _09795_/S hold703/X sky130_fd_sc_hd__mux2_1
Xhold1002 hold1002/X _15482_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 hold1024/X _15008_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 hold1057/X _15099_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ VPWR VGND VGND VPWR _08745_/Y _09694_/B _09799_/A sky130_fd_sc_hd__nor2_4
Xhold1035 hold1035/X _15297_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 hold1046/X _15295_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 hold1079/X _15302_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 hold1068/X _14887_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08676_ VPWR VGND VPWR VGND hold890/X _08562_/A _08676_/X _08691_/B1 _08675_/X _08688_/C1
+ sky130_fd_sc_hd__a221o_1
X_07627_ VPWR VGND VPWR VGND _15094_/Q _07881_/A2 _07627_/X _10074_/A0 _07159_/A _07626_/Y
+ sky130_fd_sc_hd__a221o_1
X_07558_ VPWR VGND VGND VPWR _07558_/Y _07558_/B _07558_/A sky130_fd_sc_hd__nor2_4
XFILLER_70_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07489_ VPWR VGND VGND VPWR _08603_/B _07489_/A _07489_/B sky130_fd_sc_hd__or2_1
XFILLER_10_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09228_ VGND VPWR VPWR VGND _14865_/D hold1003/X _09228_/S _09228_/A0 sky130_fd_sc_hd__mux2_1
X_13188__305 VPWR VGND VPWR VGND _14463_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_09159_ VGND VPWR VPWR VGND _14939_/D _09689_/A0 _09160_/S hold832/X sky130_fd_sc_hd__mux2_1
X_12170_ VGND VPWR VPWR VGND _12170_/X _14203_/Q _12171_/S hold230/A sky130_fd_sc_hd__mux2_1
X_11121_ VGND VPWR VPWR VGND _11121_/X hold564/A _11142_/S hold348/A sky130_fd_sc_hd__mux2_1
Xhold880 hold880/X hold880/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 hold891/X hold891/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13229__346 VPWR VGND VPWR VGND _14504_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_11052_ VPWR VGND VPWR VGND _11051_/X _11181_/A1 _11050_/X _11052_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_1044 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_77_846 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10003_ VGND VPWR _10007_/B _15617_/Q _15616_/Q _10003_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_27_1077 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14811_ _14811_/Q clkload19/A _14811_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11954_ VGND VPWR VPWR VGND _11954_/X hold766/A _11954_/S hold849/A sky130_fd_sc_hd__mux2_1
X_14742_ hold284/A _14742_/CLK _14742_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11885_ VGND VPWR VGND VPWR _11885_/X _12164_/A _11880_/X _11884_/X _12184_/C1 sky130_fd_sc_hd__o211a_1
X_14673_ hold397/A _14673_/CLK _14673_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10905_ VGND VPWR VPWR VGND _10909_/B _14790_/Q _10919_/S _14241_/Q sky130_fd_sc_hd__mux2_1
X_10836_ VGND VPWR VGND VPWR _10836_/X hold970/A _11215_/A2 _10835_/X _11205_/A sky130_fd_sc_hd__o211a_1
X_10767_ VGND VPWR VPWR VGND _10767_/X hold947/A _11091_/S hold684/A sky130_fd_sc_hd__mux2_1
XFILLER_41_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10698_ VPWR VGND VPWR VGND _10695_/X _10698_/A1 _10697_/X _10698_/X sky130_fd_sc_hd__a21o_1
X_12506_ VGND VPWR VGND VPWR _12506_/X _12670_/A1 _12502_/X _12505_/X _12670_/C1 sky130_fd_sc_hd__o211a_1
X_15225_ hold222/A _15225_/CLK _15225_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12437_ VGND VPWR VPWR VGND _12437_/X hold774/A _12661_/S hold991/A sky130_fd_sc_hd__mux2_1
X_15156_ _15156_/Q _15156_/CLK _15156_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12368_ VPWR VGND VPWR VGND _12367_/X _12376_/B2 _12366_/X _12368_/X sky130_fd_sc_hd__a21o_1
X_11319_ VPWR VGND _14825_/D _11319_/B _11327_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_12299_ VGND VPWR VGND VPWR _12299_/X _15018_/Q _12746_/A2 _11810_/S _12298_/X sky130_fd_sc_hd__o211a_1
X_15087_ _15087_/Q clkload50/A _15087_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_41_1019 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08530_ VPWR VGND VPWR VGND _08534_/B1 hold1436/X _08503_/A _08531_/B hold1401/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13022__139 VPWR VGND VPWR VGND _14265_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_08461_ VGND VPWR VGND VPWR _08461_/X hold1302/X _08458_/B _08460_/X _08919_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_36_776 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07412_ VPWR VGND VGND VPWR _07410_/Y _08287_/B _07984_/S _07412_/X sky130_fd_sc_hd__o21a_1
X_08392_ VGND VPWR VPWR VGND _15385_/D fanout41/X _08393_/S hold568/X sky130_fd_sc_hd__mux2_1
X_13373__490 VPWR VGND VPWR VGND _14648_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_07343_ VPWR VGND VPWR VGND _07665_/A _07653_/A _07403_/A _07343_/X sky130_fd_sc_hd__a21o_1
X_07274_ VGND VPWR VGND VPWR _07270_/Y _08041_/B _07981_/B _07273_/X sky130_fd_sc_hd__a21oi_2
X_09013_ VPWR VGND VGND VPWR _09890_/A _09013_/B _09013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_1424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold154 hold154/X hold154/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/X hold176/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/X hold165/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13720__837 VPWR VGND VPWR VGND _15060_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_09915_ VPWR VGND VPWR VGND _09914_/Y _09916_/B _09917_/A _14139_/D sky130_fd_sc_hd__a21oi_1
Xfanout612 VPWR VGND _07954_/S _08251_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout623 _09798_/S _09790_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold187 hold187/X hold187/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 hold198/X hold198/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 VPWR VGND _08772_/S _08745_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_09846_ VGND VPWR VPWR VGND _14176_/D hold405/X _09864_/S fanout48/X sky130_fd_sc_hd__mux2_1
Xfanout634 VPWR VGND _09675_/S _09690_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout656 _09482_/S _09451_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout667 VPWR VGND _09213_/S _09228_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout645 VGND VPWR _09521_/X _09553_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout689 VPWR VGND _08318_/S _08335_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout678 _09094_/S _09092_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09777_ VGND VPWR VPWR VGND _14272_/D _07890_/X _09795_/S hold999/X sky130_fd_sc_hd__mux2_1
XFILLER_46_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08728_ VPWR VGND VPWR VGND hold1462/X _08523_/B _08728_/X _08728_/B1 _14380_/Q _08730_/B1
+ sky130_fd_sc_hd__a221o_1
X_13614__731 VPWR VGND VPWR VGND _14954_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_08659_ VPWR VGND VPWR VGND _08664_/B _07110_/Y _08667_/A2 _08659_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11670_ VGND VPWR VGND VPWR _11670_/X hold809/A _12118_/A2 _12180_/S _11669_/X sky130_fd_sc_hd__o211a_1
XFILLER_41_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_1302 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_74_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10621_ VGND VPWR VPWR VGND _10621_/X hold801/A _10627_/S hold430/A sky130_fd_sc_hd__mux2_1
X_10552_ VGND VPWR VPWR VGND _10552_/X hold995/A _10554_/S hold899/A sky130_fd_sc_hd__mux2_1
XFILLER_10_654 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14196__914 _14196_/D _14196__914/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_1081 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10483_ VGND VPWR VPWR VGND _10483_/X hold794/A _10484_/B hold788/A sky130_fd_sc_hd__mux2_1
X_12222_ VGND VPWR VGND VPWR _12222_/X _12230_/C1 _12221_/X _12218_/X _12222_/C1 sky130_fd_sc_hd__o211a_1
X_15010_ _15010_/Q _15010_/CLK _15010_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_78_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12153_ VPWR VGND VGND VPWR _12153_/X hold241/A _12155_/S sky130_fd_sc_hd__or2_1
X_11104_ VPWR VGND VPWR VGND _11103_/X _10333_/A _11104_/B1 _11104_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12084_ VPWR VGND VPWR VGND _12083_/X _12473_/A _12491_/B1 _12084_/X sky130_fd_sc_hd__a21o_1
XFILLER_42_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11035_ VPWR VGND VGND VPWR _11035_/X hold358/A _11251_/B sky130_fd_sc_hd__or2_1
XFILLER_45_573 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14725_ hold708/A _14725_/CLK _14725_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13357__474 VPWR VGND VPWR VGND _14632_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_11937_ VPWR VGND VGND VPWR _11918_/Y _11936_/X _10562_/B _15454_/Q _15454_/D _11937_/C1
+ sky130_fd_sc_hd__o221a_1
X_14656_ hold379/A _14656_/CLK _14656_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11868_ VPWR VGND VGND VPWR _11868_/X hold161/A _12171_/S sky130_fd_sc_hd__or2_1
X_11799_ VGND VPWR VPWR VGND _11799_/X _14257_/Q _12589_/S hold152/A sky130_fd_sc_hd__mux2_1
X_10819_ VPWR VGND _10819_/X _10809_/X _10805_/X _11218_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
X_14587_ hold442/A _14587_/CLK _14587_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15208_ hold181/A _15208_/CLK _15208_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15139_ _15139_/Q _15139_/CLK _15139_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07961_ VPWR VGND VGND VPWR _15560_/Q _07990_/A _07962_/B sky130_fd_sc_hd__nor2_1
X_09700_ VGND VPWR VPWR VGND _14343_/D fanout78/X _09710_/S hold564/X sky130_fd_sc_hd__mux2_1
X_07892_ VPWR VGND VGND VPWR _15352_/Q _07892_/Y clone13/A sky130_fd_sc_hd__nand2_1
X_09631_ VGND VPWR VPWR VGND _14439_/D hold941/X _09637_/S fanout78/X sky130_fd_sc_hd__mux2_1
X_09562_ VGND VPWR VPWR VGND _14503_/D hold751/X _09584_/S fanout78/X sky130_fd_sc_hd__mux2_1
X_08513_ VPWR VGND VPWR VGND _08534_/B1 hold1421/X _08503_/A _08514_/B _15329_/Q sky130_fd_sc_hd__a22o_1
XFILLER_36_540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09493_ VGND VPWR VPWR VGND _14566_/D _09514_/S clone47/X hold1221/X sky130_fd_sc_hd__mux2_4
XFILLER_58_1368 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08444_ VPWR VGND VGND VPWR _08444_/X _15354_/Q _08488_/B sky130_fd_sc_hd__or2_1
XFILLER_51_598 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08375_ VGND VPWR VPWR VGND _15398_/D hold517/X _08375_/S fanout95/X sky130_fd_sc_hd__mux2_1
XFILLER_23_289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07326_ VGND VPWR _07325_/Y _07416_/A _07326_/Y _07154_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_17_1054 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07257_ VPWR VGND VGND VPWR _07272_/D _15458_/Q _07258_/B sky130_fd_sc_hd__or2_1
X_12957__74 VPWR VGND VPWR VGND _14200_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_13150__267 VPWR VGND VPWR VGND _14425_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_07188_ VPWR VGND _07188_/X _07189_/B _15456_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_65_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout420 VGND VPWR fanout424/X _11185_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout431 VPWR VGND _10745_/C1 _10505_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout453 VGND VPWR _07593_/X _12869_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout464 VGND VPWR _12118_/A2 _12192_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout442 VGND VPWR _10507_/A _10618_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout475 VGND VPWR _12094_/S _12086_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout497 VPWR VGND fanout497/X _07568_/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_59_676 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout486 VPWR VGND _12005_/S fanout497/X VPWR VGND sky130_fd_sc_hd__buf_2
X_09829_ VGND VPWR VPWR VGND _14223_/D _09829_/A1 _09830_/S hold347/X sky130_fd_sc_hd__mux2_1
X_12840_ VPWR VGND VGND VPWR _12842_/B _12840_/Y _12840_/B sky130_fd_sc_hd__nand2_1
X_13044__161 VPWR VGND VPWR VGND _14287_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_12771_ VGND VPWR VGND VPWR _15550_/Q _12768_/X _12770_/X _15550_/D _12807_/B1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_510 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14510_ hold275/A _14510_/CLK _14510_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11722_ VGND VPWR VPWR VGND _11722_/X _11719_/X _12396_/S _11718_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15490_ hold750/A _15490_/CLK _15490_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11653_ VGND VPWR VPWR VGND _11653_/X hold681/A _11954_/S hold297/A sky130_fd_sc_hd__mux2_1
X_14441_ hold934/A _14441_/CLK _14441_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout71 VGND VPWR _07673_/X fanout71/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_14372_ hold955/A _14372_/CLK _14372_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout60 VPWR VGND fanout60/X _07700_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_10604_ VGND VPWR VPWR VGND _10604_/X _14553_/Q _10604_/S hold245/A sky130_fd_sc_hd__mux2_1
Xfanout82 VPWR VGND VGND VPWR clone45/A clone49/A sky130_fd_sc_hd__buf_8
Xfanout93 VGND VPWR fanout94/X fanout93/X VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_11584_ VGND VPWR VPWR VGND _11585_/B _11583_/Y _12102_/S _11575_/Y sky130_fd_sc_hd__mux2_1
X_10535_ VGND VPWR VPWR VGND _10535_/X _14199_/Q _10700_/S hold324/A sky130_fd_sc_hd__mux2_1
XFILLER_10_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10466_ VGND VPWR VGND VPWR _10466_/X _10486_/A1 _10462_/X _10465_/X _10704_/C1 sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_23_Left_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12205_ VGND VPWR VPWR VGND _12209_/B hold749/A _12205_/S hold334/A sky130_fd_sc_hd__mux2_1
XFILLER_69_407 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10397_ VGND VPWR VPWR VGND _10397_/X hold933/A _10702_/S hold686/A sky130_fd_sc_hd__mux2_1
X_12136_ VGND VPWR VGND VPWR _12136_/X _12156_/A1 _12132_/X _12135_/X _12202_/C1 sky130_fd_sc_hd__o211a_1
X_12067_ VGND VPWR VPWR VGND _12067_/X hold898/A _12219_/S hold799/A sky130_fd_sc_hd__mux2_1
X_11018_ VGND VPWR VPWR VGND _11018_/X _14212_/Q _11165_/S hold205/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Left_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14708_ hold674/A _14708_/CLK _14708_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14639_ hold429/A _14639_/CLK _14639_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08160_ VPWR VGND VPWR VGND _08180_/C _08180_/B _08180_/A _08181_/A sky130_fd_sc_hd__a21o_1
XFILLER_14_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07111_ VPWR VGND VPWR VGND _09954_/B _14126_/Q sky130_fd_sc_hd__inv_2
X_08091_ VGND VPWR VGND VPWR _08091_/X _08299_/A2 _15617_/Q _08075_/X _08090_/Y sky130_fd_sc_hd__a211o_2
XPHY_EDGE_ROW_41_Left_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkload30 VGND VPWR VPWR VGND clkload30/A clkload30/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload52 clkload52/Y clkload52/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload41 VGND VPWR VPWR VGND clkload41/A clkload41/Y sky130_fd_sc_hd__clkinv_2
X_08993_ VGND VPWR VGND VPWR _08993_/X _09873_/A _09016_/B1 hold904/X _08992_/Y sky130_fd_sc_hd__a211o_1
X_13028__145 VPWR VGND VPWR VGND _14271_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07944_ VGND VPWR VGND VPWR _07944_/X _07966_/A _10066_/C _07941_/Y _10071_/A sky130_fd_sc_hd__o211a_1
X_13791__908 VPWR VGND VPWR VGND _15163_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07875_ _07876_/B _07311_/B _07897_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_25_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09614_ VGND VPWR VPWR VGND _14454_/D fanout12/X _09625_/S hold631/X sky130_fd_sc_hd__mux2_1
X_13832__949 VPWR VGND VPWR VGND _15204_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_09545_ VGND VPWR VPWR VGND _14517_/D fanout9/A _09553_/S hold180/X sky130_fd_sc_hd__mux2_1
XFILLER_52_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09476_ VGND VPWR VPWR VGND _14580_/D fanout6/X _09478_/S hold330/X sky130_fd_sc_hd__mux2_1
X_08427_ VGND VPWR VGND VPWR _08427_/X hold1282/X _08485_/A2 _08426_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
X_13685__802 VPWR VGND VPWR VGND _15025_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_36_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkload2 VGND VPWR VPWR VGND clkload2/A clkload2/Y sky130_fd_sc_hd__clkinvlp_4
X_08358_ VGND VPWR VPWR VGND _15415_/D hold591/X _08366_/S fanout37/X sky130_fd_sc_hd__mux2_1
X_13726__843 VPWR VGND VPWR VGND _15098_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_08289_ VPWR VGND VGND VPWR _15584_/Q _08289_/B _08289_/Y sky130_fd_sc_hd__nor2_1
X_07309_ VPWR VGND VPWR VGND _07811_/B _07309_/C _07811_/A _07313_/A sky130_fd_sc_hd__or3_1
X_10320_ VGND VPWR VGND VPWR _10320_/X _11259_/C1 _10315_/X _10319_/X _10765_/S sky130_fd_sc_hd__o211a_1
X_10251_ VGND VPWR VPWR VGND _10251_/X hold832/A _10258_/B hold578/A sky130_fd_sc_hd__mux2_1
XFILLER_79_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10182_ VGND VPWR VPWR VGND _10182_/X _15001_/Q _10479_/S hold777/A sky130_fd_sc_hd__mux2_1
Xfanout250 VPWR VGND _12596_/C1 _12666_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
X_14990_ hold471/A _14990_/CLK _14990_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout261 VGND VPWR _12213_/S _12694_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout272 VGND VPWR _10583_/A2 _10629_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout283 VGND VPWR _10609_/S _10602_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_75_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout294 VPWR VGND _10520_/S fanout314/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_75_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12823_ VPWR VGND _12823_/X _12821_/X _12820_/Y _12822_/A _09975_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_15611_ _15611_/Q clkload27/A _15611_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_46_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12754_ VPWR VGND VPWR VGND _12752_/Y _15545_/Q _12807_/B1 _15545_/D _12753_/X sky130_fd_sc_hd__a22o_1
XFILLER_15_532 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15542_ hold294/A _15542_/CLK _15542_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14072__1189 VPWR VGND VPWR VGND _15491_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_43_874 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11705_ VGND VPWR VPWR VGND _11705_/X hold719/A _12716_/S hold290/A sky130_fd_sc_hd__mux2_1
X_12685_ VPWR VGND VPWR VGND _12684_/X _12703_/A1 _12683_/X _12685_/Y sky130_fd_sc_hd__a21oi_1
X_15473_ _15473_/Q clkload40/A _15473_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11636_ VPWR VGND VGND VPWR _11636_/X hold549/A _12089_/S sky130_fd_sc_hd__or2_1
X_14424_ hold898/A _14424_/CLK _14424_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11567_ VGND VPWR _15444_/D _15444_/Q _11567_/A _11567_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14355_ hold861/A _14355_/CLK _14355_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xmax_cap406 VGND VPWR _07872_/Y fanout405/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold709 hold709/X hold709/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14286_ hold259/A _14286_/CLK _14286_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13469__586 VPWR VGND VPWR VGND _14744_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_10518_ VGND VPWR VGND VPWR _10518_/X hold669/A _10633_/A2 _10517_/X _10288_/S sky130_fd_sc_hd__o211a_1
X_11498_ VGND VPWR VPWR VGND _15083_/D _11497_/X _11538_/S _15083_/Q sky130_fd_sc_hd__mux2_1
XFILLER_13_1282 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10449_ VPWR VGND _10449_/X _10439_/X _10435_/X _10737_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
X_12119_ VGND VPWR VGND VPWR _12119_/X _12116_/X _12118_/X _12119_/A1 _12193_/C1 sky130_fd_sc_hd__a211o_1
Xhold1409 _09131_/A _14966_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07660_ VGND VPWR VPWR VGND _15540_/D _07954_/S clone111/X hold1197/X sky130_fd_sc_hd__mux2_4
X_07591_ VPWR VGND VPWR VGND _07591_/Y _07591_/A sky130_fd_sc_hd__inv_2
XFILLER_0_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09330_ VGND VPWR VPWR VGND _14714_/D hold723/X _09336_/S fanout29/X sky130_fd_sc_hd__mux2_1
XFILLER_34_896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09261_ VGND VPWR VPWR VGND _14782_/D fanout23/X _09275_/S hold384/X sky130_fd_sc_hd__mux2_1
X_13413__530 VPWR VGND VPWR VGND _14688_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_08212_ VGND VPWR VGND VPWR _08198_/X _10058_/A1 _08211_/X _08212_/X _08209_/X sky130_fd_sc_hd__a211o_4
X_09192_ VGND VPWR VPWR VGND _14899_/D hold362/X _09197_/S _09550_/A1 sky130_fd_sc_hd__mux2_1
X_08143_ _08143_/X _08140_/X _08141_/X _08142_/X _08294_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08074_ VGND VPWR VPWR VGND _08074_/X _08072_/X _08197_/S _07645_/X sky130_fd_sc_hd__mux2_1
X_12927__44 VPWR VGND VPWR VGND _14170_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
XFILLER_31_1382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_66_1423 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08976_ VGND VPWR VGND VPWR _15112_/D hold758/X _08985_/A2 _08975_/X _08955_/A sky130_fd_sc_hd__o211a_1
X_13262__379 VPWR VGND VPWR VGND _14537_/CLK clkload54/A sky130_fd_sc_hd__inv_2
XFILLER_29_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07927_ VPWR VGND VPWR VGND _15084_/Q _10072_/B _07927_/X _10074_/A0 _07286_/B _07926_/Y
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_1394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07858_ VGND VPWR VGND VPWR _07858_/X _07857_/A _12831_/B _07857_/Y _10071_/A sky130_fd_sc_hd__o211a_1
XFILLER_44_605 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07789_ VPWR VGND VPWR VGND _07736_/B _15556_/Q _07788_/X _07790_/B sky130_fd_sc_hd__a21o_1
X_09528_ VGND VPWR VPWR VGND _14534_/D _09537_/S fanout72/X hold1139/X sky130_fd_sc_hd__mux2_4
XFILLER_25_841 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09459_ VGND VPWR VPWR VGND _14597_/D fanout70/X _09467_/S hold389/X sky130_fd_sc_hd__mux2_1
X_13156__273 VPWR VGND VPWR VGND _14431_/CLK clkload51/A sky130_fd_sc_hd__inv_2
XFILLER_40_877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12470_ VGND VPWR VPWR VGND _12470_/X _12467_/X _12470_/S _12466_/X sky130_fd_sc_hd__mux2_1
X_11421_ VPWR VGND VPWR VGND _11421_/B _11421_/D _11421_/C _11421_/A _11421_/X sky130_fd_sc_hd__or4_2
XFILLER_61_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11352_ VGND VPWR VPWR VGND _14839_/D _14930_/Q _11355_/S hold1175/X sky130_fd_sc_hd__mux2_1
X_14140_ _14140_/Q _14140_/CLK _14140_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10303_ VPWR VGND VPWR VGND _10302_/X _10507_/A _12047_/B1 _10303_/X sky130_fd_sc_hd__a21o_1
X_11283_ VGND VPWR _11408_/A _11341_/A _14800_/D _11539_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_4_789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10234_ VGND VPWR VPWR VGND _10234_/X hold804/A _10258_/B hold461/A sky130_fd_sc_hd__mux2_1
X_10165_ VGND VPWR VPWR VGND _10165_/X _14189_/Q _10464_/S hold201/A sky130_fd_sc_hd__mux2_1
XFILLER_48_955 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14973_ hold759/A _14973_/CLK _14973_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10096_ VGND VPWR VGND VPWR _10096_/X _10614_/A1 _10092_/X _10095_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
X_13854__971 VPWR VGND VPWR VGND _15226_/CLK clkload33/A sky130_fd_sc_hd__inv_2
XFILLER_75_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12806_ VPWR VGND VGND VPWR _12817_/A _12806_/Y _12806_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_690 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10998_ VPWR VGND VGND VPWR _10998_/X hold179/A _11231_/S sky130_fd_sc_hd__or2_1
XFILLER_42_170 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12737_ VGND VPWR VGND VPWR _12737_/X _14966_/Q _12743_/A2 _12737_/B1 _12736_/X sky130_fd_sc_hd__o211a_1
X_15525_ hold352/A _15525_/CLK _15525_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15456_ _15456_/Q clkload11/A _15456_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12668_ VPWR VGND VGND VPWR _12668_/X hold208/A _12671_/S sky130_fd_sc_hd__or2_1
X_11619_ VGND VPWR VPWR VGND _11619_/X _11616_/X _12100_/S _11615_/X sky130_fd_sc_hd__mux2_1
X_14407_ _14407_/Q clkload34/A _14407_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_15387_ _15387_/Q _15387_/CLK _15387_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12599_ VGND VPWR VPWR VGND _12599_/X _15393_/Q _12599_/S _15540_/Q sky130_fd_sc_hd__mux2_1
XFILLER_15_1366 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold506 hold506/X hold506/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 hold517/X hold517/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14338_ hold713/A _14338_/CLK _14338_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold539 hold539/X hold539/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ hold908/A _14269_/CLK _14269_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold528 hold528/X hold528/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08830_ VGND VPWR VPWR VGND _15183_/D fanout44/X _08844_/S hold501/X sky130_fd_sc_hd__mux2_1
Xhold1206 hold1206/X _14135_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 hold1217/X _15336_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 hold1228/X _14147_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 hold1239/X _15151_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ VGND VPWR VPWR VGND _15245_/D fanout39/X _08776_/S hold182/X sky130_fd_sc_hd__mux2_1
XFILLER_39_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13099__216 VPWR VGND VPWR VGND _14342_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07712_ VPWR VGND VGND VPWR _07803_/A _15563_/Q _07713_/B sky130_fd_sc_hd__or2_1
X_08692_ VGND VPWR VGND VPWR _15284_/D hold1008/X _08701_/A2 _08691_/X _11937_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07643_ VPWR VGND VPWR VGND _07643_/B _07643_/C _07643_/A _07643_/X sky130_fd_sc_hd__or3_4
XFILLER_0_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07574_ VPWR VGND VGND VPWR _08214_/A _07574_/A _08232_/B sky130_fd_sc_hd__nand2_2
X_09313_ VPWR VGND VGND VPWR hold1357/X _09327_/S _09313_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09244_ _14799_/D fanout91/X fanout87/X _09242_/Y _09243_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_60_clk clkload16/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_33_1433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09175_ VGND VPWR VPWR VGND _14916_/D _09191_/S hold1147/X fanout54/X sky130_fd_sc_hd__mux2_4
X_08126_ VGND VPWR _08126_/B _12776_/A _08126_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_08057_ VGND VPWR _08058_/B _08057_/A _08057_/B VPWR VGND sky130_fd_sc_hd__xnor2_2
X_13797__914 VPWR VGND VPWR VGND _15169_/CLK clkload55/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13838__955 VPWR VGND VPWR VGND _15210_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_14071__1188 VPWR VGND VPWR VGND _15490_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_08959_ VGND VPWR VPWR VGND _08960_/B _07549_/B _09906_/A hold588/A sky130_fd_sc_hd__mux2_1
X_11970_ VGND VPWR VPWR VGND _11970_/X _11969_/X _12139_/S _11961_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10921_ VGND VPWR VPWR VGND _10921_/X _10920_/X _11244_/S _10919_/X sky130_fd_sc_hd__mux2_1
X_10852_ VGND VPWR VGND VPWR _10852_/X _11112_/A _10848_/X _10851_/X _11259_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_77_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10783_ VPWR VGND _10783_/X _10782_/X _10778_/X _10765_/S _10774_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_38_1355 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15310_ hold990/A _15310_/CLK _15310_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12522_ VGND VPWR VGND VPWR _12522_/X _12519_/X _12521_/X _12737_/B1 _12739_/C1 sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_51_clk _12972__89/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_15241_ hold593/A _15241_/CLK _15241_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12453_ VPWR VGND _12453_/X _12452_/X _12448_/X _12694_/S _12444_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11404_ VGND VPWR _11362_/X _14855_/Q _11404_/Y _11408_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_15172_ hold812/A _15172_/CLK _15172_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12384_ VGND VPWR VPWR VGND _12384_/X _14337_/Q _12408_/S _15249_/Q sky130_fd_sc_hd__mux2_1
X_11335_ VPWR VGND VPWR VGND _14829_/Q _14830_/Q _14831_/Q _11336_/B sky130_fd_sc_hd__a21oi_1
X_11266_ VPWR VGND VGND VPWR _11247_/Y _11265_/X _12751_/A2 _14410_/Q _14410_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
X_10217_ VGND VPWR VPWR VGND _10217_/X _14865_/Q _10972_/S hold530/A sky130_fd_sc_hd__mux2_1
XFILLER_80_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11197_ VPWR VGND VGND VPWR _11197_/X _11213_/S _11197_/B sky130_fd_sc_hd__or2_1
X_10148_ VGND VPWR VGND VPWR _10148_/X _15482_/Q _10633_/A2 _10147_/X _10625_/S sky130_fd_sc_hd__o211a_1
X_14956_ _14956_/Q _14956_/CLK _14956_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10079_ VGND VPWR VGND VPWR _12833_/B _12833_/A _10079_/X sky130_fd_sc_hd__or2_4
XFILLER_48_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13590__707 VPWR VGND VPWR VGND _14921_/CLK clkload48/A sky130_fd_sc_hd__inv_2
XFILLER_63_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14887_ _14887_/Q _14887_/CLK _14887_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13631__748 VPWR VGND VPWR VGND _14971_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_15508_ _15508_/Q _15508_/CLK _15508_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_clk clkload50/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07290_ VPWR VGND VGND VPWR _14402_/Q _07301_/A2 _07301_/B1 _07292_/B sky130_fd_sc_hd__o21a_1
X_15439_ _15439_/Q clkload47/A _15439_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13484__601 VPWR VGND VPWR VGND _14759_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
XFILLER_50_1076 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold325 hold325/X hold325/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 hold314/X hold314/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 hold303/X hold303/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13525__642 VPWR VGND VPWR VGND _14805_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_09931_ VPWR VGND VGND VPWR _09931_/C _09931_/B _14134_/Q _09931_/Y sky130_fd_sc_hd__nor3_1
Xhold358 hold358/X hold358/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 hold336/X hold336/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 hold347/X hold347/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 hold369/X hold369/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout805 VPWR VGND _11382_/S fanout829/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout816 VGND VPWR fanout829/X _12233_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout838 VPWR VGND _08943_/A _11567_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout827 VGND VPWR _11347_/A _08571_/B VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_63_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout849 VPWR VGND _07668_/B _07422_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_09862_ VGND VPWR VPWR VGND _14160_/D hold395/X _09867_/S _09862_/A0 sky130_fd_sc_hd__mux2_1
Xhold1014 _09878_/A _14150_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ VGND VPWR VPWR VGND _15196_/D fanout98/X _08814_/S hold186/X sky130_fd_sc_hd__mux2_1
X_09793_ VGND VPWR VPWR VGND _14256_/D _09862_/A0 _09798_/S hold394/X sky130_fd_sc_hd__mux2_1
Xhold1003 hold1003/X _14865_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 hold1058/X _15100_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ VPWR VGND VPWR VGND _09311_/B _09694_/B _09240_/A _09556_/C sky130_fd_sc_hd__or3b_2
XFILLER_39_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1025 hold1025/X _15292_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 hold1036/X _15278_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 hold1047/X _15028_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 hold1069/X _15006_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_744 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08675_ VGND VPWR VPWR VGND _08675_/X _14400_/Q _08684_/S _14384_/Q sky130_fd_sc_hd__mux2_1
XFILLER_54_788 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07626_ VPWR VGND VGND VPWR _07626_/A _07972_/B _07626_/Y sky130_fd_sc_hd__nor2_1
X_07557_ VGND VPWR VGND VPWR _07555_/B _07557_/X _07560_/B _07557_/D _07555_/A sky130_fd_sc_hd__and4bb_2
Xclkbuf_leaf_33_clk clkload51/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07488_ _07489_/B _07486_/C _07486_/B _07486_/A _07487_/A _08608_/B VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__o311a_1
X_09227_ VGND VPWR VPWR VGND _14866_/D hold993/X _09228_/S _09829_/A1 sky130_fd_sc_hd__mux2_1
X_09158_ VGND VPWR VPWR VGND _14940_/D _09550_/A1 _09163_/S hold856/X sky130_fd_sc_hd__mux2_1
X_08109_ VGND VPWR VPWR VGND _15523_/D fanout10/X _08267_/S hold248/X sky130_fd_sc_hd__mux2_1
X_09089_ VGND VPWR VPWR VGND _15004_/D hold1101/X _09094_/S _09688_/A0 sky130_fd_sc_hd__mux2_1
X_11120_ VGND VPWR VPWR VGND _11120_/X hold751/A _11142_/S hold643/A sky130_fd_sc_hd__mux2_1
Xhold881 hold881/X hold881/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13268__385 VPWR VGND VPWR VGND _14543_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
Xhold870 hold870/X hold870/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ VGND VPWR VPWR VGND _11051_/X _11048_/X _11162_/S _11047_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold892 hold892/X hold892/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10002_ VGND VPWR VPWR VGND _10002_/A _15616_/D _10003_/C sky130_fd_sc_hd__xor2_1
X_14810_ _14810_/Q _14810_/CLK _14810_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14741_ hold304/A _14741_/CLK _14741_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11953_ VGND VPWR VGND VPWR _11953_/X _12189_/C1 _11948_/X _11952_/X _12139_/S sky130_fd_sc_hd__o211a_1
X_11884_ VPWR VGND VGND VPWR _11884_/X _11958_/A _11884_/B sky130_fd_sc_hd__or2_1
X_14672_ hold671/A _14672_/CLK _14672_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10904_ VPWR VGND VPWR VGND _10903_/X _10930_/C1 _10902_/X _10904_/Y sky130_fd_sc_hd__a21oi_1
X_10835_ VPWR VGND VGND VPWR _10835_/X hold246/A _10835_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_24_clk clkload31/A clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_10766_ VPWR VGND VGND VPWR _11173_/A _10766_/B _10766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_1016 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_9_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10697_ VPWR VGND VPWR VGND _10696_/X _10677_/S _10697_/B1 _10697_/X sky130_fd_sc_hd__a21o_1
X_12505_ VPWR VGND VGND VPWR _12505_/X _12536_/S _12505_/B sky130_fd_sc_hd__or2_1
XFILLER_9_689 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15224_ hold171/A _15224_/CLK _15224_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12436_ VPWR VGND VGND VPWR _12658_/A _12436_/B _12436_/Y sky130_fd_sc_hd__nor2_1
X_15155_ _15155_/Q _15155_/CLK _15155_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13509__626 VPWR VGND VPWR VGND _14784_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
XFILLER_12_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12367_ VGND VPWR VPWR VGND _12367_/X _12364_/X _12367_/S _12363_/X sky130_fd_sc_hd__mux2_1
X_11318_ VGND VPWR VPWR VGND _11319_/B _11317_/X _14825_/Q _11313_/C sky130_fd_sc_hd__mux2_1
X_12298_ VPWR VGND VGND VPWR _12298_/X hold891/A _12708_/S sky130_fd_sc_hd__or2_1
X_15086_ _15086_/Q clkload50/A _15086_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_79_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11249_ VGND VPWR VPWR VGND _11249_/X _14378_/Q _11251_/B _14730_/Q sky130_fd_sc_hd__mux2_1
X_13899__1016 VPWR VGND VPWR VGND _15271_/CLK clkload27/A sky130_fd_sc_hd__inv_2
XFILLER_48_571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13061__178 VPWR VGND VPWR VGND _14304_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_14939_ hold832/A _14939_/CLK _14939_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08460_ VPWR VGND VGND VPWR _08460_/X _15346_/Q _08486_/B sky130_fd_sc_hd__or2_1
X_08391_ VGND VPWR VPWR VGND _15386_/D fanout45/X _08405_/S hold826/X sky130_fd_sc_hd__mux2_1
X_07411_ VPWR VGND VGND VPWR _07411_/A _10074_/S _08287_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_15_clk clkload23/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07342_ VPWR VGND VPWR VGND _07652_/A _07653_/A _07340_/X _07403_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_950 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14070__1187 VPWR VGND VPWR VGND _15489_/CLK clkload19/A sky130_fd_sc_hd__inv_2
XFILLER_32_994 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07273_ VGND VPWR VGND VPWR _07273_/X _07268_/A _07272_/X _07264_/B _07262_/X sky130_fd_sc_hd__a211o_1
X_09012_ VGND VPWR VGND VPWR _15100_/D hold1058/X _09015_/A2 _09011_/X _11327_/A sky130_fd_sc_hd__o211a_1
Xhold177 hold177/X hold177/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/X hold166/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/X hold155/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ VGND VPWR _09931_/B hold1152/X _09914_/Y _14140_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xfanout602 _08773_/S _08776_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold188 hold188/X hold188/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 VGND VPWR _07132_/Y _08251_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold199 hold199/X hold199/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout624 VPWR VGND _09790_/S _09764_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout635 VGND VPWR _09660_/X _09690_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout657 VPWR VGND _09345_/S _09336_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout646 VPWR VGND _09549_/S _09552_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09845_ VGND VPWR VPWR VGND _14177_/D hold628/X _09864_/S clone5/X sky130_fd_sc_hd__mux2_1
X_13302__419 VPWR VGND VPWR VGND _14577_/CLK clkload51/A sky130_fd_sc_hd__inv_2
Xfanout668 _09228_/S _09198_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout679 VGND VPWR _09061_/X _09092_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_46_508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09776_ VGND VPWR VPWR VGND _14273_/D _09792_/S fanout52/X hold1251/X sky130_fd_sc_hd__mux2_4
X_08727_ VGND VPWR VGND VPWR _15270_/D hold977/X _08731_/A2 _08726_/X _11294_/A sky130_fd_sc_hd__o211a_1
X_13653__770 VPWR VGND VPWR VGND _14993_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_08658_ VGND VPWR VGND VPWR _15294_/D hold1034/X _08704_/A2 _08657_/X _08717_/C1
+ sky130_fd_sc_hd__o211a_1
X_07609_ VGND VPWR VGND VPWR _07609_/X _07857_/A _07606_/X _07608_/Y _10071_/A sky130_fd_sc_hd__o211a_1
XFILLER_74_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08589_ VGND VPWR VGND VPWR _08589_/X _08617_/A _08627_/C1 hold865/X _08588_/Y sky130_fd_sc_hd__a211o_1
XFILLER_74_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10620_ VGND VPWR VGND VPWR _10620_/X _14876_/Q _10633_/A2 _10619_/X _10625_/S sky130_fd_sc_hd__o211a_1
X_10551_ VGND VPWR VPWR VGND _10555_/B hold417/A _10554_/S hold402/A sky130_fd_sc_hd__mux2_1
X_10482_ VGND VPWR VGND VPWR _10482_/X _10479_/X _10481_/X _10486_/A1 _10697_/B1 sky130_fd_sc_hd__a211o_1
X_12221_ VGND VPWR VPWR VGND _12221_/X _12220_/X _12221_/S _12219_/X sky130_fd_sc_hd__mux2_1
X_12152_ VGND VPWR VGND VPWR _12152_/X _12149_/X _12151_/X _12156_/A1 _12212_/A1 sky130_fd_sc_hd__a211o_1
X_11103_ VGND VPWR VPWR VGND _11103_/X _14889_/Q _11109_/S _15425_/Q sky130_fd_sc_hd__mux2_1
XFILLER_46_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12083_ VPWR VGND _12083_/X _12082_/X _12078_/X _12213_/S _12074_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_46_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11034_ VGND VPWR VPWR VGND _11034_/X hold775/A _11251_/B hold527/A sky130_fd_sc_hd__mux2_1
XFILLER_49_346 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14724_ hold561/A _14724_/CLK _14724_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11936_ VPWR VGND VPWR VGND _11935_/X _12214_/A _11973_/B _11936_/X sky130_fd_sc_hd__a21o_1
X_14655_ hold741/A _14655_/CLK _14655_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11867_ VGND VPWR VGND VPWR _11867_/X _11864_/X _11866_/X _11958_/A _12175_/A1 sky130_fd_sc_hd__a211o_1
X_11798_ VGND VPWR VPWR VGND _11802_/B hold605/A _12589_/S hold308/A sky130_fd_sc_hd__mux2_1
XFILLER_53_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10818_ VPWR VGND VGND VPWR _10815_/X _10817_/X _10765_/S _10818_/X sky130_fd_sc_hd__o21a_1
X_14586_ hold218/A _14586_/CLK _14586_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_13_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10749_ VGND VPWR VPWR VGND _10753_/B hold619/A _11091_/S hold376/A sky130_fd_sc_hd__mux2_1
X_15207_ hold324/A _15207_/CLK _15207_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_57_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12419_ VGND VPWR VPWR VGND _12423_/B hold567/A _12661_/S hold559/A sky130_fd_sc_hd__mux2_1
X_15138_ _15138_/Q _15138_/CLK _15138_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07960_ VPWR VGND VPWR VGND _08002_/B1 _15623_/Q _08002_/A2 _07960_/X _15587_/Q sky130_fd_sc_hd__a22o_1
X_15069_ _15069_/Q clkload15/A _15069_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_4_clk _12951__68/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_13596__713 VPWR VGND VPWR VGND _14936_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_07891_ VGND VPWR VPWR VGND _07954_/S fanout49/X hold1109/X _15534_/D sky130_fd_sc_hd__mux2_2
XFILLER_60_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09630_ VGND VPWR VPWR VGND _09637_/S hold1203/X fanout81/X _14440_/D sky130_fd_sc_hd__mux2_2
X_13637__754 VPWR VGND VPWR VGND _14977_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_3_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09561_ VGND VPWR VPWR VGND _09584_/S hold1165/X clone49/X _14504_/D sky130_fd_sc_hd__mux2_2
X_08512_ VPWR VGND _15330_/D _08512_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_71_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09492_ VGND VPWR VPWR VGND _14567_/D fanout79/X _09514_/S hold456/X sky130_fd_sc_hd__mux2_1
X_08443_ VGND VPWR VGND VPWR _15355_/D _15354_/Q _08448_/B _08442_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
X_08374_ VGND VPWR VPWR VGND _15399_/D hold345/X _08375_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
X_07325_ VPWR VGND VGND VPWR _07612_/A _07606_/B _07325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07256_ VPWR VGND VGND VPWR _14392_/Q _07230_/S _07265_/B1 _07258_/B sky130_fd_sc_hd__o21a_1
X_07187_ VPWR VGND VGND VPWR _14390_/Q _07230_/S _07265_/B1 _07189_/B sky130_fd_sc_hd__o21a_1
X_12972__89 VPWR VGND VPWR VGND _14215_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
XFILLER_79_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout421 VGND VPWR _11104_/B1 _11259_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout432 VGND VPWR _07851_/Y _10505_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout410 VGND VPWR _10704_/C1 _10697_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout465 VPWR VGND _12118_/A2 _12080_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout443 VGND VPWR _10729_/A _10507_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout454 VPWR VGND _10617_/S _10469_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout487 VGND VPWR _11882_/S _12171_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_47_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09828_ VGND VPWR VPWR VGND _14224_/D _09862_/A0 _09833_/S hold229/X sky130_fd_sc_hd__mux2_1
Xfanout476 VGND VPWR _11628_/S _12094_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout498 VGND VPWR _12205_/S _12155_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_73_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09759_ VGND VPWR VPWR VGND _14287_/D _09829_/A1 _09760_/S hold255/X sky130_fd_sc_hd__mux2_1
X_12770_ VPWR VGND _12770_/X _12788_/S _08155_/X _12789_/A _12769_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_70_842 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_42_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11721_ VGND VPWR VGND VPWR _11721_/X _12720_/A1 _11717_/X _11720_/X _12720_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_14_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_758 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11652_ VGND VPWR VPWR VGND _11652_/X _14189_/Q _11954_/S hold201/A sky130_fd_sc_hd__mux2_1
X_14204__922 _14204_/D _14204__922/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_14440_ _14440_/Q _14440_/CLK _14440_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout50 VPWR VGND fanout50/X _07890_/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout72 VPWR VGND fanout72/X _07659_/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout83 VPWR VGND VGND VPWR fanout86/X fanout83/X sky130_fd_sc_hd__buf_8
X_13430__547 VPWR VGND VPWR VGND _14705_/CLK clkload54/A sky130_fd_sc_hd__inv_2
Xfanout61 VPWR VGND VPWR VGND fanout61/X _07700_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10603_ VGND VPWR VPWR VGND _10603_/X hold451/A _10612_/S hold593/A sky130_fd_sc_hd__mux2_1
X_14371_ hold776/A _14371_/CLK _14371_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13898__1015 VPWR VGND VPWR VGND _15270_/CLK clkload27/A sky130_fd_sc_hd__inv_2
Xfanout94 VPWR VGND fanout94/X _07424_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_11583_ VPWR VGND VPWR VGND _11582_/X _12101_/A1 _11581_/X _11583_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10534_ VGND VPWR VGND VPWR _10534_/X _10634_/C1 _10529_/X _10533_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
X_10465_ VPWR VGND VGND VPWR _10465_/X _10467_/S _10465_/B sky130_fd_sc_hd__or2_1
X_13283__400 VPWR VGND VPWR VGND _14558_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_10396_ VPWR VGND VGND VPWR _10507_/A _10396_/B _10396_/Y sky130_fd_sc_hd__nor2_1
X_12204_ VPWR VGND VPWR VGND _12203_/X _12212_/A1 _12202_/X _12204_/Y sky130_fd_sc_hd__a21oi_1
X_12135_ VPWR VGND VGND VPWR _12135_/X _12147_/S _12135_/B sky130_fd_sc_hd__or2_1
X_13324__441 VPWR VGND VPWR VGND _14599_/CLK clkload42/A sky130_fd_sc_hd__inv_2
XFILLER_1_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12066_ VPWR VGND VGND VPWR _12473_/A _12066_/B _12066_/Y sky130_fd_sc_hd__nor2_1
X_11017_ VGND VPWR VPWR VGND _11017_/X hold392/A _11054_/S hold370/A sky130_fd_sc_hd__mux2_1
XFILLER_77_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14707_ hold710/A _14707_/CLK _14707_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_33_544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11919_ VPWR VGND VGND VPWR _11919_/X hold612/A _12149_/S sky130_fd_sc_hd__or2_1
XFILLER_33_566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14638_ hold635/A _14638_/CLK _14638_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07110_ VPWR VGND VPWR VGND _07110_/Y _14380_/Q sky130_fd_sc_hd__inv_2
X_14569_ hold415/A _14569_/CLK _14569_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08090_ VGND VPWR _08088_/X _08089_/X _08090_/Y _10059_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
Xclkload20 VGND VPWR VGND VPWR clkload20/Y clkload20/A sky130_fd_sc_hd__inv_12
Xclkload31 VPWR VGND VGND VPWR clkload31/Y clkload31/A sky130_fd_sc_hd__inv_16
Xclkload53 VPWR VGND VPWR VGND clkload53/Y clkload53/A sky130_fd_sc_hd__inv_6
Xclkload42 VPWR VGND VGND VPWR clkload42/Y clkload42/A sky130_fd_sc_hd__inv_16
X_08992_ VPWR VGND VGND VPWR _09873_/A _08992_/B _08992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_1384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13067__184 VPWR VGND VPWR VGND _14310_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_07943_ VPWR VGND _10066_/C _07943_/B _07943_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07874_ VPWR VGND VPWR VGND _10890_/A _08286_/A clone17/X _07890_/C sky130_fd_sc_hd__a21oi_1
X_09613_ VGND VPWR VPWR VGND _14455_/D fanout16/X _09625_/S hold1005/X sky130_fd_sc_hd__mux2_1
X_13871__988 VPWR VGND VPWR VGND _15243_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_09544_ VGND VPWR VPWR VGND _14518_/D fanout14/X _09555_/S hold236/X sky130_fd_sc_hd__mux2_1
X_09475_ VGND VPWR VPWR VGND _14581_/D fanout9/X _09485_/S hold497/X sky130_fd_sc_hd__mux2_1
X_08426_ VPWR VGND VGND VPWR _08426_/X _15363_/Q _08484_/B sky130_fd_sc_hd__or2_1
XFILLER_36_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08357_ VGND VPWR VPWR VGND _15416_/D hold452/X _08372_/S fanout39/X sky130_fd_sc_hd__mux2_1
Xclkload3 VGND VPWR VPWR VGND clkload3/A clkload3/Y sky130_fd_sc_hd__clkinvlp_4
X_13765__882 VPWR VGND VPWR VGND _15137_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_08288_ _08289_/B _07418_/B _15582_/Q _10075_/B _08286_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07308_ VPWR VGND VPWR VGND _07859_/A _07899_/A _07876_/A _07820_/A _07309_/C sky130_fd_sc_hd__or4_1
XFILLER_50_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07239_ VGND VPWR VGND VPWR _08156_/B _08162_/A _08135_/B _07206_/X sky130_fd_sc_hd__a21oi_2
X_10250_ VGND VPWR VGND VPWR _10250_/X hold993/A _11003_/A2 _10249_/X _10911_/S sky130_fd_sc_hd__o211a_1
X_13308__425 VPWR VGND VPWR VGND _14583_/CLK clkload9/A sky130_fd_sc_hd__inv_2
XFILLER_78_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10181_ VGND VPWR VPWR VGND _10185_/B hold984/A _10479_/S hold653/A sky130_fd_sc_hd__mux2_1
Xfanout240 VGND VPWR _08270_/A1 _12212_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout251 VPWR VGND _12666_/A1 _07955_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout262 VPWR VGND _12472_/S _12213_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout273 VGND VPWR _10583_/A2 _10688_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_43_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout295 VGND VPWR _10472_/S _10687_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout284 VGND VPWR _10140_/S _10609_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_47_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15610_ _15610_/Q clkload27/A _15610_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_75_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_74_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12822_ VPWR VGND VGND VPWR _12822_/A _12822_/B _12822_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_894 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12753_ VPWR VGND VGND VPWR _10079_/X _07769_/A _08257_/X _12789_/A _12753_/X _12807_/A1
+ sky130_fd_sc_hd__o221a_1
X_15541_ hold164/A _15541_/CLK _15541_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15472_ _15472_/Q clkload51/A _15472_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11704_ VGND VPWR VGND VPWR _11704_/X _12722_/A1 _11699_/X _11703_/X _12864_/A1 sky130_fd_sc_hd__o211a_1
X_12684_ VGND VPWR VPWR VGND _12684_/X _12681_/X _12684_/S _12680_/X sky130_fd_sc_hd__mux2_1
X_14423_ hold887/A _14423_/CLK _14423_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11635_ VGND VPWR VPWR VGND _11635_/X hold498/A _12089_/S hold727/A sky130_fd_sc_hd__mux2_1
X_11566_ VPWR VGND VPWR VGND _11565_/Y _11567_/C _11542_/A _15443_/D sky130_fd_sc_hd__a21oi_1
X_14354_ hold965/A _14354_/CLK _14354_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14285_ hold278/A _14285_/CLK _14285_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10517_ VPWR VGND VGND VPWR _10517_/X hold236/A _10521_/B sky130_fd_sc_hd__or2_1
X_11497_ VGND VPWR VPWR VGND _11497_/X _11496_/X _11537_/S _15463_/Q sky130_fd_sc_hd__mux2_1
X_10448_ VPWR VGND VGND VPWR _10445_/X _10447_/X clone2/X _10448_/X sky130_fd_sc_hd__o21a_1
X_10379_ VGND VPWR VPWR VGND _10383_/B hold806/A _10390_/S hold443/A sky130_fd_sc_hd__mux2_1
X_12118_ VGND VPWR VGND VPWR _12118_/X _15013_/Q _12118_/A2 _12118_/B1 _12117_/X sky130_fd_sc_hd__o211a_1
X_12049_ VGND VPWR VPWR VGND _12053_/B hold760/A _12219_/S hold654/A sky130_fd_sc_hd__mux2_1
XFILLER_26_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_19_850 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07590_ VPWR VGND VPWR VGND clone20/A _15160_/Q _07589_/X _07591_/A sky130_fd_sc_hd__a21oi_1
X_13101__218 VPWR VGND VPWR VGND _14344_/CLK clkload41/A sky130_fd_sc_hd__inv_2
XFILLER_34_875 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09260_ VGND VPWR VPWR VGND _14783_/D fanout27/X _09268_/S hold721/X sky130_fd_sc_hd__mux2_1
X_08211_ VGND VPWR VGND VPWR _08206_/X _08147_/A _08210_/Y _08211_/X _08249_/B2 sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13749__866 VPWR VGND VPWR VGND _15121_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_09191_ VGND VPWR VPWR VGND _14900_/D hold353/X _09191_/S _09653_/A0 sky130_fd_sc_hd__mux2_1
X_08142_ VGND VPWR VGND VPWR _08280_/A2 _07204_/B _08104_/B _08142_/X _08137_/A sky130_fd_sc_hd__a2bb2o_1
X_08073_ VPWR VGND VGND VPWR _11440_/B _08197_/S _08073_/B sky130_fd_sc_hd__nand2_1
X_13969__1086 VPWR VGND VPWR VGND _15341_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_12942__59 VPWR VGND VPWR VGND _14185_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_08975_ VGND VPWR VGND VPWR _08975_/X _08983_/A _08972_/A hold1445/X _08974_/Y sky130_fd_sc_hd__a211o_1
XFILLER_75_208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07926_ VPWR VGND VGND VPWR _07926_/A _07972_/B _07926_/Y sky130_fd_sc_hd__nor2_1
X_07857_ VPWR VGND VGND VPWR _07857_/A _07857_/Y _07857_/B sky130_fd_sc_hd__nand2_1
X_13897__1014 VPWR VGND VPWR VGND _15269_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_07788_ _07788_/X _08037_/B _08037_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_56_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_44_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09527_ VGND VPWR VPWR VGND _14535_/D fanout77/X _09549_/S hold421/X sky130_fd_sc_hd__mux2_1
XFILLER_80_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09458_ VGND VPWR VPWR VGND _14598_/D _09467_/S fanout74/X hold1120/X sky130_fd_sc_hd__mux2_4
XFILLER_61_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08409_ VGND VPWR VPWR VGND _15368_/D _09691_/A0 _08409_/S hold426/X sky130_fd_sc_hd__mux2_1
X_09389_ VGND VPWR VPWR VGND _14660_/D hold592/X _09408_/S fanout65/X sky130_fd_sc_hd__mux2_1
X_11420_ VGND VPWR VPWR VGND _11420_/X _14820_/Q _11420_/S hold1166/X sky130_fd_sc_hd__mux2_1
X_11351_ VGND VPWR VPWR VGND _14838_/D _14929_/Q _11355_/S hold1262/X sky130_fd_sc_hd__mux2_1
XFILLER_3_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10302_ VPWR VGND _10302_/X _10301_/X _10297_/X _10617_/S _10293_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11282_ VGND VPWR VGND VPWR _11567_/C _15444_/Q _11410_/A sky130_fd_sc_hd__or2_4
XFILLER_3_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_3_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10233_ VGND VPWR VPWR VGND _10233_/X hold664/A _10258_/B hold267/A sky130_fd_sc_hd__mux2_1
X_13542__659 VPWR VGND VPWR VGND _14873_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_10164_ VGND VPWR VGND VPWR _10164_/X _10693_/B1 _10159_/X _10163_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
X_10095_ VPWR VGND VGND VPWR _10095_/X _10613_/A _10095_/B sky130_fd_sc_hd__or2_1
X_14972_ hold433/A _14972_/CLK _14972_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13395__512 VPWR VGND VPWR VGND _14670_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XFILLER_47_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12805_ VPWR VGND VGND VPWR _12822_/A _12805_/Y _12805_/B sky130_fd_sc_hd__nand2_1
X_13436__553 VPWR VGND VPWR VGND _14711_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_15524_ hold216/A _15524_/CLK _15524_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10997_ VGND VPWR VPWR VGND _10997_/X hold810/A _11231_/S hold204/A sky130_fd_sc_hd__mux2_1
X_12736_ VPWR VGND VGND VPWR _12736_/X _14925_/Q _12736_/B sky130_fd_sc_hd__or2_1
X_15455_ _15455_/Q clkload32/A _15455_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12667_ VGND VPWR VPWR VGND _12667_/X hold657/A _12671_/S hold294/A sky130_fd_sc_hd__mux2_1
X_15386_ hold826/A _15386_/CLK _15386_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14406_ _14406_/Q clkload49/A _14406_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11618_ VGND VPWR VGND VPWR _11618_/X _11638_/A1 _11614_/X _11617_/X _12115_/C1 sky130_fd_sc_hd__o211a_1
X_12598_ VGND VPWR VGND VPWR _12598_/X _15508_/Q _12746_/A2 _12367_/S _12597_/X sky130_fd_sc_hd__o211a_1
X_14337_ _14337_/Q _14337_/CLK _14337_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_580 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11549_ VPWR VGND VGND VPWR _11549_/A _11549_/Y _11549_/B sky130_fd_sc_hd__nand2_1
Xhold518 hold518/X hold518/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 hold507/X hold507/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 hold529/X hold529/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ hold544/A _14268_/CLK _14268_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14199_ _14199_/Q _14199_/CLK _14199_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1207 hold1207/X _14497_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1218 _15337_/D _08479_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ VGND VPWR VPWR VGND _15246_/D clone44/A _08773_/S hold321/X sky130_fd_sc_hd__mux2_1
Xhold1229 hold1229/X _14494_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07711_ VGND VPWR VPWR VGND _07713_/B _15590_/Q _07807_/S _07519_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_978 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14092__1209 VPWR VGND VPWR VGND _15511_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_08691_ VPWR VGND VPWR VGND hold1465/X _08700_/A2 _08691_/X _08691_/B1 _08690_/X
+ _08700_/B1 sky130_fd_sc_hd__a221o_1
X_07642_ _07643_/C _07638_/X _07639_/Y _07641_/X _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09312_ VPWR VGND VPWR VGND _09312_/X _09729_/A _09660_/B sky130_fd_sc_hd__or2_2
X_07573_ VPWR VGND VGND VPWR _07573_/A _08233_/B _07573_/B sky130_fd_sc_hd__nand2_1
X_13179__296 VPWR VGND VPWR VGND _14454_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
XFILLER_34_683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_61_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09243_ VPWR VGND VGND VPWR _09243_/X _09243_/A _09269_/S sky130_fd_sc_hd__or2_1
XFILLER_22_878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_33_1445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09174_ VGND VPWR VPWR VGND _14917_/D hold834/X _09191_/S clone55/X sky130_fd_sc_hd__mux2_1
X_08125_ VGND VPWR VPWR VGND _08128_/B _08124_/X _08099_/B _12833_/A _08299_/A2 _15615_/Q
+ sky130_fd_sc_hd__a32o_1
X_08056_ _08057_/B _07738_/X _08056_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_13877__994 VPWR VGND VPWR VGND _15249_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_08958_ VGND VPWR VGND VPWR _15118_/D hold988/X _08985_/A2 _08957_/X _08955_/A sky130_fd_sc_hd__o211a_1
X_08889_ VGND VPWR VGND VPWR _15148_/D hold1179/X _08893_/A2 _08888_/X _11974_/C1
+ sky130_fd_sc_hd__o211a_1
X_07909_ VGND VPWR VPWR VGND _07909_/A _12821_/A _07909_/B sky130_fd_sc_hd__xor2_1
X_13123__240 VPWR VGND VPWR VGND _14366_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_10920_ VGND VPWR VPWR VGND _10920_/X hold843/A _11146_/B hold465/A sky130_fd_sc_hd__mux2_1
X_10851_ VPWR VGND VGND VPWR _10851_/X _10851_/A _10851_/B sky130_fd_sc_hd__or2_1
X_10782_ VGND VPWR VGND VPWR _10782_/X _10781_/X _10780_/X _11215_/C1 _11217_/C1 sky130_fd_sc_hd__a211o_1
X_12521_ VGND VPWR VGND VPWR _12521_/X hold914/A _12669_/A2 _12735_/S _12520_/X sky130_fd_sc_hd__o211a_1
X_15240_ hold220/A _15240_/CLK _15240_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_8_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12452_ VGND VPWR VGND VPWR _12452_/X _12451_/X _12450_/X _12662_/A1 _12662_/C1 sky130_fd_sc_hd__a211o_1
X_11403_ VGND VPWR VPWR VGND _14854_/D _11402_/X _11401_/Y _11396_/X _11395_/X _14854_/Q
+ sky130_fd_sc_hd__a32o_1
X_15171_ hold399/A _15171_/CLK _15171_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12383_ VGND VPWR VPWR VGND _12383_/X _14497_/Q _12408_/S hold628/A sky130_fd_sc_hd__mux2_1
X_11334_ VGND VPWR _11338_/B _14830_/Q _14831_/Q _14829_/Q VPWR VGND sky130_fd_sc_hd__and3_1
X_11265_ VPWR VGND VPWR VGND _11264_/X _11247_/A _12750_/B1 _11265_/X sky130_fd_sc_hd__a21o_1
X_12987__104 VPWR VGND VPWR VGND _14230_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_14039__1156 VPWR VGND VPWR VGND _15411_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_10216_ VGND VPWR VGND VPWR _10216_/X hold967/A _11003_/A2 _10215_/X _11004_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_80_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11196_ VGND VPWR VPWR VGND _11196_/X hold415/A _11204_/S hold234/A sky130_fd_sc_hd__mux2_1
X_10147_ VPWR VGND VGND VPWR _10147_/X hold250/A _10632_/B sky130_fd_sc_hd__or2_1
X_14955_ hold817/A _14955_/CLK _14955_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10078_ VPWR VGND VGND VPWR _10078_/A _12833_/B _10078_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_63_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07129__1 VPWR VGND VPWR VGND _14126_/CLK clkload25/A sky130_fd_sc_hd__inv_2
XFILLER_63_734 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14886_ hold964/A _14886_/CLK _14886_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13968__1085 VPWR VGND VPWR VGND _15340_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_13670__787 VPWR VGND VPWR VGND _15010_/CLK clkload6/A sky130_fd_sc_hd__inv_2
Xclkbuf_0_clk VGND VPWR VGND VPWR clk clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_15507_ _15507_/Q _15507_/CLK _15507_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12719_ VPWR VGND VGND VPWR _12719_/X _12721_/S _12719_/B sky130_fd_sc_hd__or2_1
X_15438_ _15438_/Q clkload47/A _15438_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13896__1013 VPWR VGND VPWR VGND _15268_/CLK clkload20/A sky130_fd_sc_hd__inv_2
XFILLER_11_1017 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15369_ hold719/A _15369_/CLK _15369_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold304 hold304/X hold304/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 hold315/X hold315/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 hold326/X hold326/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ VGND VPWR VPWR VGND _14134_/D hold1359/X _09931_/B _09929_/X sky130_fd_sc_hd__mux2_1
Xhold359 hold359/X hold359/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 hold337/X hold337/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 hold348/X hold348/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13564__681 VPWR VGND VPWR VGND _14895_/CLK clkload7/A sky130_fd_sc_hd__inv_2
Xfanout806 VPWR VGND _08925_/C1 fanout829/X VPWR VGND sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout839 VGND VPWR _07544_/B _11567_/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout828 VGND VPWR fanout829/X _08571_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09861_ VGND VPWR VPWR VGND _14161_/D hold551/X _09861_/S _08190_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout817 VPWR VGND _11388_/S _11974_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
X_12912__29 VPWR VGND VPWR VGND _14155_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_08812_ VGND VPWR VPWR VGND _15197_/D _09865_/A0 _08814_/S hold201/X sky130_fd_sc_hd__mux2_1
Xhold1015 hold1015/X _14485_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ VGND VPWR VPWR VGND _14257_/D _09792_/A1 _09792_/S hold1065/X sky130_fd_sc_hd__mux2_1
Xhold1004 hold1004/X _15009_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13107__224 VPWR VGND VPWR VGND _14350_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
Xhold1048 _09875_/A _14151_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ VPWR VGND _15259_/D _08743_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
Xhold1026 hold1026/X _14878_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1037 hold1037/X _14437_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 hold1059/X _15281_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08674_ VGND VPWR VGND VPWR _15290_/D hold1127/X _08701_/A2 _08673_/X _12085_/C1
+ sky130_fd_sc_hd__o211a_1
X_07625_ VPWR VGND VGND VPWR _07625_/A _10075_/A _07625_/Y sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07556_ VGND VPWR _07557_/D _07556_/B _08956_/B _07560_/D VPWR VGND sky130_fd_sc_hd__and3_1
X_07487_ VPWR VGND VGND VPWR _07487_/A _08609_/A _07487_/B sky130_fd_sc_hd__nand2_1
X_09226_ VGND VPWR VPWR VGND _14867_/D hold778/X _09231_/S _09550_/A1 sky130_fd_sc_hd__mux2_1
XFILLER_10_859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09157_ VGND VPWR VPWR VGND _14941_/D _09653_/A0 _09157_/S hold975/X sky130_fd_sc_hd__mux2_1
X_13805__922 VPWR VGND VPWR VGND _15177_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_08108_ VGND VPWR VGND VPWR _08108_/X _08099_/Y _08107_/X _12833_/A _08095_/X sky130_fd_sc_hd__a211o_1
X_09088_ VGND VPWR VPWR VGND _15005_/D hold1033/X _09088_/S _09792_/A1 sky130_fd_sc_hd__mux2_1
X_08039_ VGND VPWR VPWR VGND _08039_/X _08038_/X _07837_/Y _12833_/A _08037_/Y _07810_/A
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold882 hold882/X hold882/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold860 hold860/X hold860/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 hold871/X hold871/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold893 hold893/X hold893/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ VGND VPWR VGND VPWR _11050_/X _11185_/A1 _11046_/X _11049_/X _11185_/C1 sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_10_Left_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10001_ VPWR VGND VGND VPWR _10003_/C _10001_/B _15615_/D sky130_fd_sc_hd__nor2_1
XFILLER_79_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14740_ hold312/A _14740_/CLK _14740_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11952_ VGND VPWR VGND VPWR _11952_/X _11949_/X _11951_/X _11968_/S _12185_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_45_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11883_ VGND VPWR VPWR VGND _11883_/X hold910/A _12183_/S hold725/A sky130_fd_sc_hd__mux2_1
X_10903_ VGND VPWR VPWR VGND _10903_/X _10900_/X _10911_/S _10899_/X sky130_fd_sc_hd__mux2_1
X_14671_ hold638/A _14671_/CLK _14671_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10834_ VGND VPWR VPWR VGND _10834_/X hold706/A _10835_/B hold244/A sky130_fd_sc_hd__mux2_1
X_10765_ VGND VPWR VPWR VGND _10766_/B _10764_/Y _10765_/S _10756_/Y sky130_fd_sc_hd__mux2_1
XFILLER_40_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12504_ VGND VPWR VPWR VGND _12504_/X hold587/A _12652_/S hold441/A sky130_fd_sc_hd__mux2_1
X_12978__95 VPWR VGND VPWR VGND _14221_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_10696_ VGND VPWR VPWR VGND _10696_/X _14878_/Q _10696_/S hold380/A sky130_fd_sc_hd__mux2_1
XFILLER_9_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15223_ _15223_/Q _15223_/CLK _15223_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12435_ VGND VPWR VPWR VGND _12436_/B _12434_/Y _12731_/S _12426_/Y sky130_fd_sc_hd__mux2_1
X_14091__1208 VPWR VGND VPWR VGND _15510_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_12366_ VGND VPWR VGND VPWR _12366_/X _12367_/S _12361_/X _12365_/X _12863_/A1 sky130_fd_sc_hd__o211a_1
X_15154_ _15154_/Q _15154_/CLK _15154_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13548__665 VPWR VGND VPWR VGND _14879_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_11317_ VGND VPWR VGND VPWR _11317_/X _11421_/B _14833_/Q _11316_/Y sky130_fd_sc_hd__a21bo_1
X_12297_ VGND VPWR VPWR VGND _12297_/X hold853/A _12708_/S hold663/A sky130_fd_sc_hd__mux2_1
X_15085_ _15085_/Q clkload50/A _15085_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11248_ VGND VPWR VPWR VGND _11248_/X _14442_/Q _11251_/B _14698_/Q sky130_fd_sc_hd__mux2_1
XFILLER_80_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11179_ VGND VPWR VPWR VGND _11179_/X _14891_/Q _11179_/S hold448/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14938_ hold967/A _14938_/CLK _14938_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14869_ hold827/A _14869_/CLK _14869_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08390_ VGND VPWR VPWR VGND _08393_/S fanout49/X hold1178/X _15387_/D sky130_fd_sc_hd__mux2_2
X_07410_ VPWR VGND VGND VPWR _07410_/C _07410_/B _07416_/A _07410_/Y sky130_fd_sc_hd__nor3_1
X_07341_ _07652_/A _07319_/B _15471_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_07272_ VGND VPWR _07272_/C _08010_/A _07272_/X _07272_/D _08025_/A VPWR VGND sky130_fd_sc_hd__and4b_1
X_09011_ VGND VPWR VGND VPWR _09011_/X _09890_/A _09016_/B1 hold1057/X _09010_/Y sky130_fd_sc_hd__a211o_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold156 hold156/X hold156/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/X hold167/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ VPWR VGND VPWR VGND _14139_/Q _09931_/B _14140_/Q _09916_/B sky130_fd_sc_hd__or3_1
Xfanout603 _08776_/S _08745_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold189 hold189/X hold189/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 hold178/X hold178/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 VGND VPWR _11480_/S _11477_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout625 _09792_/S _09795_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout647 VPWR VGND _09537_/S _09552_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout636 _09625_/S _09617_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09844_ VGND VPWR VPWR VGND _14178_/D hold825/X _09861_/S fanout57/X sky130_fd_sc_hd__mux2_1
Xfanout658 VPWR VGND _09336_/S _09312_/X VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_74_807 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout669 VPWR VGND _09197_/S _09188_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_13341__458 VPWR VGND VPWR VGND _14616_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
XFILLER_39_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09775_ VGND VPWR VPWR VGND _14274_/D fanout58/X _09792_/S hold552/X sky130_fd_sc_hd__mux2_1
X_08726_ VPWR VGND VPWR VGND _15269_/Q _09912_/A _08726_/X _08728_/B1 _14381_/Q _08726_/C1
+ sky130_fd_sc_hd__a221o_1
X_08657_ VPWR VGND VPWR VGND hold1452/X _08714_/A2 _08657_/X _08711_/B1 _08656_/X
+ _08722_/C1 sky130_fd_sc_hd__a221o_1
X_13194__311 VPWR VGND VPWR VGND _14469_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_07608_ VGND VPWR _07607_/Y _07857_/A _07608_/Y _07410_/C VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_74_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08588_ VPWR VGND VGND VPWR _08617_/A _08992_/B _08588_/Y sky130_fd_sc_hd__nor2_1
X_14038__1155 VPWR VGND VPWR VGND _15410_/CLK clkload10/A sky130_fd_sc_hd__inv_2
XFILLER_74_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07539_ VPWR VGND VGND VPWR _07539_/A _07539_/B _07539_/Y _07539_/C sky130_fd_sc_hd__nand3_1
X_13235__352 VPWR VGND VPWR VGND _14510_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_10550_ VPWR VGND VPWR VGND _10547_/X _10634_/A1 _10549_/X _10550_/X sky130_fd_sc_hd__a21o_1
X_10481_ VGND VPWR VGND VPWR _10481_/X _15491_/Q _10688_/A2 _10480_/X _10467_/S sky130_fd_sc_hd__o211a_1
X_09209_ VGND VPWR VPWR VGND _14884_/D hold966/X _09213_/S clone5/X sky130_fd_sc_hd__mux2_1
X_12220_ VGND VPWR VPWR VGND _12220_/X hold913/A _12220_/S hold418/A sky130_fd_sc_hd__mux2_1
X_13967__1084 VPWR VGND VPWR VGND _15339_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_12151_ VGND VPWR VGND VPWR _12151_/X _15014_/Q _12229_/A2 _12147_/S _12150_/X sky130_fd_sc_hd__o211a_1
XFILLER_78_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11102_ VGND VPWR VPWR VGND _11102_/X hold458/A _11102_/S hold354/A sky130_fd_sc_hd__mux2_1
Xhold690 hold690/X hold690/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12082_ VGND VPWR VGND VPWR _12082_/X _12081_/X _12080_/X _12230_/A1 _12226_/C1 sky130_fd_sc_hd__a211o_1
X_11033_ VGND VPWR VGND VPWR _11033_/X _11181_/A1 _11032_/X _11029_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_65_807 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13895__1012 VPWR VGND VPWR VGND _15267_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
Xhold1390 _10000_/A _15615_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14723_ hold446/A _14723_/CLK _14723_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11935_ VPWR VGND _11935_/X _11934_/X _11930_/X _12139_/S _11926_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14654_ _14654_/Q _14654_/CLK _14654_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_27_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11866_ VGND VPWR VGND VPWR _11866_/X _14483_/Q _12192_/A2 _12174_/S _11865_/X sky130_fd_sc_hd__o211a_1
X_11797_ VPWR VGND VPWR VGND _11796_/X _12744_/C1 _11795_/X _11797_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10817_ VGND VPWR VGND VPWR _10817_/X _10851_/A _10813_/X _10816_/X _11263_/C1 sky130_fd_sc_hd__o211a_1
X_14585_ hold245/A _14585_/CLK _14585_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10748_ VPWR VGND VGND VPWR _10729_/Y _10747_/X _10562_/B _14396_/Q _14396_/D _11937_/C1
+ sky130_fd_sc_hd__o221a_1
X_13782__899 VPWR VGND VPWR VGND _15154_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_10679_ VGND VPWR VGND VPWR _10679_/X hold938/A _10688_/A2 _10678_/X _10698_/A1 sky130_fd_sc_hd__o211a_1
X_15206_ hold341/A _15206_/CLK _15206_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12418_ VPWR VGND VGND VPWR _12399_/Y _12417_/X _12751_/A2 _15467_/Q _15467_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
X_12349_ VPWR VGND VGND VPWR _12349_/X hold630/A _12370_/S sky130_fd_sc_hd__or2_1
X_15137_ _15137_/Q _15137_/CLK _15137_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15068_ _15068_/Q clkload15/A _15068_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_67_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07890_ VGND VPWR VPWR VGND _07890_/D _07890_/C _07890_/B _07890_/A _07890_/X sky130_fd_sc_hd__or4_4
X_09560_ VGND VPWR VPWR VGND _14505_/D hold903/X _09584_/S clone133/X sky130_fd_sc_hd__mux2_1
XFILLER_36_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13676__793 VPWR VGND VPWR VGND _15016_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_08511_ VPWR VGND VPWR VGND _08534_/B1 _15329_/Q _08503_/A _08512_/B hold1435/X sky130_fd_sc_hd__a22o_1
XFILLER_36_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09491_ VGND VPWR VPWR VGND _14568_/D clone45/X _09514_/S hold580/X sky130_fd_sc_hd__mux2_1
X_08442_ VPWR VGND VGND VPWR _08442_/X _15355_/Q _08488_/B sky130_fd_sc_hd__or2_1
XFILLER_36_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13219__336 VPWR VGND VPWR VGND _14494_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_1_1081 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08373_ VGND VPWR VPWR VGND _15400_/D hold445/X _08375_/S _09229_/A0 sky130_fd_sc_hd__mux2_1
X_07324_ VPWR VGND VGND VPWR _07625_/A _07619_/B _07323_/Y _07606_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_943 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07255_ VGND VPWR VGND VPWR _07249_/A _08066_/A _08041_/B _07249_/B sky130_fd_sc_hd__a21oi_4
X_07186_ VPWR VGND VPWR VGND _07981_/A _07186_/A _07186_/B sky130_fd_sc_hd__or2_2
Xfanout411 VGND VPWR _08178_/A1 _10704_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout422 VGND VPWR _11104_/B1 _11217_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout400 VPWR VGND _11252_/C1 _10846_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout455 VPWR VGND _10469_/S _10728_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout444 VGND VPWR _07691_/X _10729_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout433 VPWR VGND _11237_/A1 _10891_/C1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout466 VGND VPWR _12080_/A2 _12229_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09827_ VGND VPWR VPWR VGND _14225_/D _09827_/A1 _09827_/S hold308/X sky130_fd_sc_hd__mux2_1
Xfanout488 VGND VPWR _11882_/S _11876_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout477 VGND VPWR _11628_/S _11756_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout499 VGND VPWR _12149_/S _12205_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09758_ VGND VPWR VPWR VGND _14288_/D _09862_/A0 _09763_/S hold240/X sky130_fd_sc_hd__mux2_1
X_08709_ VGND VPWR VGND VPWR _08709_/X _08714_/A2 _08722_/C1 hold872/X _08708_/X sky130_fd_sc_hd__a211o_1
X_14090__1207 VPWR VGND VPWR VGND _15509_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XFILLER_54_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11720_ VPWR VGND VGND VPWR _11720_/X _12396_/S _11720_/B sky130_fd_sc_hd__or2_1
XFILLER_15_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09689_ VGND VPWR VPWR VGND _14351_/D hold1029/X _09690_/S _09689_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_74_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11651_ VGND VPWR VPWR VGND _11651_/X _14253_/Q _11950_/B hold278/A sky130_fd_sc_hd__mux2_1
Xfanout40 VPWR VGND fanout40/X _07953_/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_70_1014 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout73 VPWR VGND fanout73/X _07659_/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout62 VGND VPWR _07700_/X fanout62/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_11582_ VGND VPWR VPWR VGND _11582_/X _11579_/X _12098_/A _11578_/X sky130_fd_sc_hd__mux2_1
X_14370_ hold866/A _14370_/CLK _14370_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10602_ VGND VPWR VPWR VGND _10602_/X _14489_/Q _10602_/S hold351/A sky130_fd_sc_hd__mux2_1
Xfanout84 VPWR VGND VGND VPWR fanout86/X fanout84/X sky130_fd_sc_hd__buf_8
X_10533_ VGND VPWR VGND VPWR _10533_/X _10532_/X _10531_/X _10625_/S _10630_/C1 sky130_fd_sc_hd__a211o_1
Xfanout95 VGND VPWR fanout96/X fanout95/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_12948__65 VPWR VGND VPWR VGND _14191_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_7_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10464_ VGND VPWR VPWR VGND _10464_/X hold596/A _10464_/S hold304/A sky130_fd_sc_hd__mux2_1
X_10395_ VGND VPWR VPWR VGND _10396_/B _10394_/Y _10469_/S _10386_/Y sky130_fd_sc_hd__mux2_1
X_12203_ VGND VPWR VPWR VGND _12203_/X _12200_/X _12221_/S _12199_/X sky130_fd_sc_hd__mux2_1
X_13012__129 VPWR VGND VPWR VGND _14255_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_12134_ VGND VPWR VPWR VGND _12134_/X hold566/A _12155_/S hold193/A sky130_fd_sc_hd__mux2_1
X_12065_ VGND VPWR VPWR VGND _12066_/B _12064_/Y _12139_/S _12056_/Y sky130_fd_sc_hd__mux2_1
X_13363__480 VPWR VGND VPWR VGND _14638_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_11016_ VGND VPWR VPWR VGND _11020_/B hold560/A _11054_/S hold364/A sky130_fd_sc_hd__mux2_1
XFILLER_46_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13710__827 VPWR VGND VPWR VGND _15050_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_14706_ hold583/A _14706_/CLK _14706_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11918_ VPWR VGND VGND VPWR _12214_/A _11918_/B _11918_/Y sky130_fd_sc_hd__nor2_1
X_14637_ hold333/A _14637_/CLK _14637_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_33_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11849_ VGND VPWR VGND VPWR _11849_/X _14942_/Q _12040_/A2 _12099_/A1 _11848_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_707 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14568_ hold580/A _14568_/CLK _14568_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkload10 clkload10/Y clkload10/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
XFILLER_9_295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14499_ _14499_/Q _14499_/CLK _14499_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkload32 clkload32/Y clkload32/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload43 clkload43/Y clkload43/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload21 VGND VPWR VGND VPWR clkload21/A clkload21/Y sky130_fd_sc_hd__bufinv_8
Xclkload54 VGND VPWR VPWR VGND clkload54/A clkload54/Y sky130_fd_sc_hd__clkinvlp_4
X_13604__721 VPWR VGND VPWR VGND _14944_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_08991_ VGND VPWR VGND VPWR hold921/A hold920/X _09015_/A2 _08990_/X _09000_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_64_1341 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07942_ VPWR VGND VPWR VGND _07942_/B _07942_/C _07945_/A _07943_/B sky130_fd_sc_hd__or3_1
X_14037__1154 VPWR VGND VPWR VGND _15409_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_07873_ VPWR VGND VPWR VGND _07873_/B1 _15353_/Q _08495_/A2 _07873_/X _15142_/Q sky130_fd_sc_hd__a22o_1
XFILLER_56_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09612_ VGND VPWR VPWR VGND _14456_/D fanout20/X _09622_/S hold744/X sky130_fd_sc_hd__mux2_1
X_09543_ VGND VPWR VPWR VGND _14519_/D fanout17/X _09555_/S hold546/X sky130_fd_sc_hd__mux2_1
X_09474_ VGND VPWR VPWR VGND _14582_/D fanout14/X _09485_/S hold668/X sky130_fd_sc_hd__mux2_1
X_08425_ VPWR VGND VGND VPWR _08425_/X _08425_/A _09937_/A sky130_fd_sc_hd__or2_1
X_13966__1083 VPWR VGND VPWR VGND _15338_/CLK clkload28/A sky130_fd_sc_hd__inv_2
XFILLER_71_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08356_ VGND VPWR VPWR VGND _15417_/D _08356_/S hold1113/X fanout42/X sky130_fd_sc_hd__mux2_4
Xclkload4 clkload4/X clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07307_ VPWR VGND VGND VPWR _07899_/A _07311_/B _07307_/B sky130_fd_sc_hd__or2_1
XFILLER_36_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08287_ VPWR VGND VGND VPWR _10075_/B _08287_/A _08287_/B sky130_fd_sc_hd__or2_1
X_07238_ VPWR VGND VPWR VGND _08179_/B _08180_/A _07209_/X _08156_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13894__1011 VPWR VGND VPWR VGND _15266_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_07169_ VPWR VGND _07668_/A _07319_/B _15471_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_79_707 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13347__464 VPWR VGND VPWR VGND _14622_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_10180_ VPWR VGND VPWR VGND _10177_/X _10486_/A1 _10179_/X _10180_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout230 VGND VPWR fanout234/X _12739_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout241 VPWR VGND _12230_/C1 _08270_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout252 VPWR VGND _12111_/C1 _12222_/C1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout263 VPWR VGND _12213_/S _07935_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout274 VGND VPWR _10583_/A2 _10744_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout296 VGND VPWR _10472_/S _10390_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout285 VGND VPWR _10140_/S _10271_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_12821_ VPWR VGND VGND VPWR _12821_/X _12821_/A _12829_/S sky130_fd_sc_hd__or2_1
XFILLER_28_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15540_ _15540_/Q _15540_/CLK _15540_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12752_ VGND VPWR _12833_/B _08256_/X _12752_/Y _07765_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_37_1207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12683_ VGND VPWR VGND VPWR _12683_/X _12256_/S _12679_/X _12682_/X _12702_/C1 sky130_fd_sc_hd__o211a_1
X_15471_ _15471_/Q clkload39/A _15471_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11703_ VGND VPWR VGND VPWR _11703_/X _11702_/X _11701_/X _12476_/S _12485_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_42_375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14422_ _14422_/Q _14422_/CLK _14422_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11634_ VGND VPWR VGND VPWR _11634_/X _11633_/X _11632_/X _12106_/S _12017_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_50_1418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11565_ VGND VPWR _11563_/B hold1287/X _11565_/Y _15442_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_50_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14353_ hold859/A _14353_/CLK _14353_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11496_ VGND VPWR VPWR VGND _11496_/X _15084_/Q _11535_/C _15082_/Q sky130_fd_sc_hd__mux2_1
X_14284_ hold541/A _14284_/CLK _14284_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_755 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10516_ VGND VPWR VPWR VGND _10516_/X hold802/A _10516_/S hold216/A sky130_fd_sc_hd__mux2_1
X_10447_ VGND VPWR VGND VPWR _10447_/X _10662_/S _10443_/X _10446_/X _10667_/C1 sky130_fd_sc_hd__o211a_1
X_10378_ VPWR VGND VGND VPWR _10359_/Y _10377_/X _10710_/B _14386_/Q _14386_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
X_12117_ VPWR VGND VGND VPWR _12117_/X hold331/A _12117_/B sky130_fd_sc_hd__or2_1
X_12048_ VPWR VGND VGND VPWR _12029_/Y _12047_/X _10710_/B _15457_/Q _15457_/D _11294_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_59_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13140__257 VPWR VGND VPWR VGND _14415_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XFILLER_61_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08210_ VGND VPWR _08210_/B _08210_/Y _08210_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_09190_ VGND VPWR VPWR VGND _14901_/D hold411/X _09197_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_08141_ VPWR VGND VPWR VGND _08293_/A3 _15073_/Q _11440_/B _08141_/X _08115_/A sky130_fd_sc_hd__a22o_1
X_08072_ VPWR VGND VPWR VGND _08252_/A2 _15343_/Q _08253_/A2 _08072_/X _15148_/Q sky130_fd_sc_hd__a22o_1
X_13034__151 VPWR VGND VPWR VGND _14277_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_08974_ VPWR VGND VGND VPWR _08983_/A _08974_/B _08974_/Y sky130_fd_sc_hd__nor2_1
X_07925_ VPWR VGND VGND VPWR _07925_/A _10075_/A _07925_/Y sky130_fd_sc_hd__nor2_1
X_07856_ VPWR VGND VGND VPWR _07856_/A _07857_/B _07856_/B sky130_fd_sc_hd__nand2_1
X_07787_ VGND VPWR _08057_/A _08056_/B _08037_/B _07738_/X VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_44_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09526_ VGND VPWR VPWR VGND _14536_/D fanout80/X _09549_/S hold208/X sky130_fd_sc_hd__mux2_1
XFILLER_25_854 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09457_ VGND VPWR VPWR VGND _14599_/D fanout79/X _09467_/S hold326/X sky130_fd_sc_hd__mux2_1
XFILLER_80_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08408_ VGND VPWR VPWR VGND _15369_/D _09228_/A0 _08408_/S hold719/X sky130_fd_sc_hd__mux2_1
X_09388_ VGND VPWR VPWR VGND _14661_/D hold365/X _09408_/S fanout69/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08339_ VPWR VGND _09834_/A _15577_/Q _09164_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_12918__35 VPWR VGND VPWR VGND _14161_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_11350_ VGND VPWR VPWR VGND _11350_/X _14928_/Q _11355_/S hold1264/X sky130_fd_sc_hd__mux2_1
X_10301_ VGND VPWR VGND VPWR _10301_/X _10300_/X _10299_/X _10523_/A1 _10630_/C1 sky130_fd_sc_hd__a211o_1
X_11281_ VPWR VGND VGND VPWR _11408_/A _11567_/C _15444_/Q sky130_fd_sc_hd__nor2_4
X_13581__698 VPWR VGND VPWR VGND _14912_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_10232_ VGND VPWR VPWR VGND _10232_/X hold968/A _10258_/B hold731/A sky130_fd_sc_hd__mux2_1
X_10163_ VGND VPWR VGND VPWR _10163_/X _10162_/X _10161_/X _10467_/S _10697_/B1 sky130_fd_sc_hd__a211o_1
XFILLER_48_902 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10094_ VGND VPWR VPWR VGND _10094_/X hold789/A _10602_/S hold165/A sky130_fd_sc_hd__mux2_1
X_14971_ hold327/A _14971_/CLK _14971_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_56_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12804_ VGND VPWR VPWR VGND _12805_/B _07990_/X _12820_/B _07993_/B sky130_fd_sc_hd__mux2_1
X_15523_ hold248/A _15523_/CLK _15523_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13475__592 VPWR VGND VPWR VGND _14750_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_15_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_16_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10996_ VGND VPWR VGND VPWR _10996_/X _11237_/A1 _10995_/X _10992_/X _12869_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_43_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12735_ VGND VPWR VPWR VGND _12735_/X _12734_/X _12735_/S _12733_/X sky130_fd_sc_hd__mux2_1
X_14036__1153 VPWR VGND VPWR VGND _15408_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_12666_ VGND VPWR VGND VPWR _12666_/X _12666_/A1 _12665_/X _12662_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_15454_ VGND VPWR VGND VPWR _15454_/Q _15454_/D clkload17/A sky130_fd_sc_hd__dfxtp_4
X_12597_ VPWR VGND VGND VPWR _12597_/X _14534_/Q _12599_/S sky130_fd_sc_hd__or2_1
X_13018__135 VPWR VGND VPWR VGND _14261_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_15385_ hold568/A _15385_/CLK _15385_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14405_ _14405_/Q clkload39/A _14405_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11617_ VPWR VGND VGND VPWR _11617_/X _12100_/S _11617_/B sky130_fd_sc_hd__or2_1
X_11548_ VPWR VGND VPWR VGND _11547_/Y _11549_/B _11542_/A _15434_/D sky130_fd_sc_hd__a21oi_1
X_14336_ hold973/A _14336_/CLK _14336_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold508 hold508/X hold508/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13822__939 VPWR VGND VPWR VGND _15194_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_14267_ hold943/A _14267_/CLK _14267_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11479_ VGND VPWR VPWR VGND _11479_/X _11478_/X _11491_/S _15457_/Q sky130_fd_sc_hd__mux2_1
Xhold519 hold519/X hold519/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14198_ _14198_/Q _14198_/CLK _14198_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13965__1082 VPWR VGND VPWR VGND _15337_/CLK clkload28/A sky130_fd_sc_hd__inv_2
XFILLER_32_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_29_Left_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_3_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1219 hold1219/X _15184_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07710_ VPWR VGND VGND VPWR _07710_/A _07888_/A _07710_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1208 hold1208/X _14337_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08690_ VGND VPWR VPWR VGND _08690_/X _14395_/Q _08690_/S _14379_/Q sky130_fd_sc_hd__mux2_1
X_07641_ VPWR VGND VPWR VGND _15093_/Q _07881_/A2 _07641_/X _10074_/A0 _07163_/A _07640_/Y
+ sky130_fd_sc_hd__a221o_1
X_13716__833 VPWR VGND VPWR VGND _15056_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_26_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13893__1010 VPWR VGND VPWR VGND _15265_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_07572_ VPWR VGND _07572_/X _07573_/B _07573_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_09311_ VPWR VGND VGND VPWR _15581_/Q _09311_/B _09660_/B _09556_/C sky130_fd_sc_hd__nand3_1
X_09242_ VPWR VGND VPWR VGND _09242_/Y _09269_/S sky130_fd_sc_hd__inv_2
X_09173_ VGND VPWR VPWR VGND _14918_/D hold382/X _09194_/S fanout62/X sky130_fd_sc_hd__mux2_1
X_08124_ VPWR VGND VGND VPWR _08124_/X _15552_/Q _08145_/A sky130_fd_sc_hd__or2_1
XFILLER_33_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12885__2 VPWR VGND VPWR VGND _14127_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08055_ VPWR VGND VGND VPWR _08214_/B _07421_/Y _08053_/X _07421_/A _08070_/A _07996_/X
+ sky130_fd_sc_hd__o221a_1
X_08957_ VGND VPWR VGND VPWR _08957_/X _08983_/A _08969_/A hold985/X _08956_/Y sky130_fd_sc_hd__a211o_1
X_08888_ VPWR VGND VGND VPWR _08888_/X _15148_/Q _08918_/B sky130_fd_sc_hd__or2_1
X_07908_ VPWR VGND VPWR VGND _15626_/Q _07929_/A2 _07908_/X _07908_/B1 _15590_/Q _07907_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07839_ VGND VPWR _07990_/A _15558_/Q _15559_/Q _08023_/A VPWR VGND sky130_fd_sc_hd__and3_1
X_13459__576 VPWR VGND VPWR VGND _14734_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_10850_ VGND VPWR VPWR VGND _10850_/X hold826/A _10850_/S hold305/A sky130_fd_sc_hd__mux2_1
X_10781_ VGND VPWR VPWR VGND _10781_/X hold599/A _10850_/S hold206/A sky130_fd_sc_hd__mux2_1
XFILLER_40_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09509_ VGND VPWR VPWR VGND _14550_/D fanout14/X _09520_/S hold822/X sky130_fd_sc_hd__mux2_1
XFILLER_24_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13989__1106 VPWR VGND VPWR VGND _15361_/CLK clkload27/A sky130_fd_sc_hd__inv_2
X_12520_ VPWR VGND VGND VPWR _12520_/X hold295/A _12671_/S sky130_fd_sc_hd__or2_1
X_12451_ VGND VPWR VPWR VGND _12451_/X hold687/A _12623_/S hold162/A sky130_fd_sc_hd__mux2_1
X_11402_ VPWR VGND _11402_/X _14853_/Q _14851_/Q _14852_/Q _14854_/Q VGND VPWR sky130_fd_sc_hd__a31o_1
X_15170_ hold562/A _15170_/CLK _15170_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XANTENNA_90 _14385_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12382_ VGND VPWR VPWR VGND _12386_/B _14625_/Q _12408_/S hold450/A sky130_fd_sc_hd__mux2_1
X_11333_ VPWR VGND VGND VPWR _11332_/X _11421_/C _11316_/Y _14830_/Q _14830_/D _11337_/C1
+ sky130_fd_sc_hd__o221a_1
X_11264_ VPWR VGND _11264_/X _11263_/X _11259_/X _10765_/S _11255_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_4_566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10215_ VPWR VGND VGND VPWR _10215_/X hold499/A _10567_/S sky130_fd_sc_hd__or2_1
XFILLER_45_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11195_ VGND VPWR VPWR VGND _11195_/X hold513/A _11204_/S hold553/A sky130_fd_sc_hd__mux2_1
X_10146_ VGND VPWR VPWR VGND _10146_/X hold704/A _10632_/B hold233/A sky130_fd_sc_hd__mux2_1
X_13403__520 VPWR VGND VPWR VGND _14678_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_14954_ hold743/A _14954_/CLK _14954_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10077_ VPWR VGND VPWR VGND _12833_/B _10071_/X _10073_/Y _10076_/X wire858/X _15576_/Q
+ sky130_fd_sc_hd__o311a_2
XFILLER_63_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14885_ _14885_/Q _14885_/CLK _14885_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10979_ VGND VPWR VPWR VGND _10983_/B hold661/A _10994_/S hold223/A sky130_fd_sc_hd__mux2_1
X_15506_ hold914/A _15506_/CLK _15506_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12718_ VGND VPWR VPWR VGND _12718_/X _14570_/Q _12726_/S _14602_/Q sky130_fd_sc_hd__mux2_1
X_15437_ _15437_/Q clkload51/A _15437_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13252__369 VPWR VGND VPWR VGND _14527_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_12649_ VGND VPWR VPWR VGND _12653_/B hold732/A _12651_/S hold276/A sky130_fd_sc_hd__mux2_1
X_15368_ hold426/A _15368_/CLK _15368_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold305 hold305/X hold305/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15299_ _15299_/Q _15299_/CLK _15299_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14319_ hold664/A _14319_/CLK _14319_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold316 hold316/X hold316/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 hold349/X hold349/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold338/X hold338/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 hold327/X hold327/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout807 VPWR VGND _11420_/S _08529_/A VPWR VGND sky130_fd_sc_hd__buf_2
X_09860_ VGND VPWR VPWR VGND _14162_/D hold474/X _09867_/S _09860_/A0 sky130_fd_sc_hd__mux2_1
Xfanout829 VGND VPWR _14154_/Q fanout829/X VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout818 VPWR VGND _08919_/C1 _11974_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
X_13146__263 VPWR VGND VPWR VGND _14421_/CLK clkload24/A sky130_fd_sc_hd__inv_2
XFILLER_58_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09791_ VGND VPWR VPWR VGND _14258_/D _09826_/A1 _09798_/S hold529/X sky130_fd_sc_hd__mux2_1
Xhold1005 hold1005/X _14455_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08811_ VGND VPWR VPWR VGND _15198_/D _09622_/A1 _08811_/S hold190/X sky130_fd_sc_hd__mux2_1
Xhold1016 hold1016/X _14496_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ VGND VPWR VPWR VGND _08743_/B _08492_/X _07560_/X _15638_/Q _09938_/C _15259_/Q
+ sky130_fd_sc_hd__a32o_1
Xhold1027 hold1027/X _14477_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 hold1049/X _15015_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_1261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1038 hold1038/X _14359_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_38_231 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08673_ VPWR VGND VPWR VGND _15289_/Q _08562_/A _08673_/X _08691_/B1 _08672_/X _08688_/C1
+ sky130_fd_sc_hd__a221o_1
X_07624_ VGND VPWR VGND VPWR _07624_/X _07984_/S _07620_/Y _07623_/Y _10071_/A sky130_fd_sc_hd__o211a_1
XFILLER_54_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07555_ VGND VPWR VGND VPWR _07555_/B _07555_/A _08174_/A _07560_/C _07554_/D sky130_fd_sc_hd__or4bb_4
XFILLER_35_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07486_ VPWR VGND VPWR VGND _07486_/B _07486_/C _07486_/A _07487_/B sky130_fd_sc_hd__or3_1
X_09225_ VGND VPWR VPWR VGND _14868_/D hold1072/X _09228_/S _09653_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_42_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_10_805 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13844__961 VPWR VGND VPWR VGND _15216_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_09156_ VGND VPWR VPWR VGND _14942_/D _09826_/A1 _09163_/S hold1091/X sky130_fd_sc_hd__mux2_1
X_08107_ VPWR VGND VPWR VGND _15616_/Q _08249_/A2 _08107_/X _08106_/X _08294_/B1 _08098_/Y
+ sky130_fd_sc_hd__a221o_1
X_09087_ VGND VPWR VPWR VGND _15006_/D hold1069/X _09094_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_08038_ VPWR VGND VPWR VGND _08059_/B _15555_/Q _15556_/Q _08038_/X sky130_fd_sc_hd__a21o_1
Xhold861 hold861/X hold861/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 hold872/X hold872/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold850 hold850/X hold850/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ VPWR VGND VGND VPWR _10000_/A _10000_/B _10001_/B sky130_fd_sc_hd__nor2_1
Xhold883 hold883/X hold883/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 hold894/X hold894/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09989_ VGND VPWR _09993_/B _15611_/Q _15610_/Q _09989_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14035__1152 VPWR VGND VPWR VGND _15407_/CLK clkload17/A sky130_fd_sc_hd__inv_2
XFILLER_76_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11951_ VGND VPWR VGND VPWR _11951_/X hold901/A _12192_/A2 _11948_/S _11950_/X sky130_fd_sc_hd__o211a_1
XFILLER_72_565 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11882_ VGND VPWR VPWR VGND _11882_/X hold835/A _11882_/S hold344/A sky130_fd_sc_hd__mux2_1
X_10902_ VGND VPWR VGND VPWR _10902_/X _11235_/A1 _10898_/X _10901_/X _10918_/C1 sky130_fd_sc_hd__o211a_1
X_14670_ hold672/A _14670_/CLK _14670_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10833_ VGND VPWR VPWR VGND _10833_/X _10832_/X _11205_/A _10831_/X sky130_fd_sc_hd__mux2_1
X_10764_ VPWR VGND VPWR VGND _10763_/X _11218_/A1 _10762_/X _10764_/Y sky130_fd_sc_hd__a21oi_1
X_13964__1081 VPWR VGND VPWR VGND _15336_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_12503_ VGND VPWR VPWR VGND _12503_/X _14212_/Q _12652_/S hold205/A sky130_fd_sc_hd__mux2_1
X_10695_ VGND VPWR VPWR VGND _10695_/X hold992/A _10696_/S hold337/A sky130_fd_sc_hd__mux2_1
XFILLER_9_647 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15222_ _15222_/Q _15222_/CLK _15222_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12434_ VPWR VGND VPWR VGND _12433_/X _12656_/A1 _12432_/X _12434_/Y sky130_fd_sc_hd__a21oi_1
X_12365_ VPWR VGND VGND VPWR _12365_/X _12375_/S _12365_/B sky130_fd_sc_hd__or2_1
X_15153_ _15153_/Q _15153_/CLK _15153_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_66_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13089__206 VPWR VGND VPWR VGND _14332_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_11316_ VGND VPWR _11421_/C _14822_/Q _11316_/Y _11410_/A VPWR VGND sky130_fd_sc_hd__o21ai_2
X_15084_ _15084_/Q clkload15/A _15084_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12296_ VGND VPWR VGND VPWR _12296_/X _12703_/A1 _12291_/X _12295_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_80_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11247_ VPWR VGND VGND VPWR _11247_/A _11247_/B _11247_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11178_ VGND VPWR VGND VPWR _11178_/X hold813/A _11184_/A2 _11177_/X _11178_/C1 sky130_fd_sc_hd__o211a_1
X_10129_ VGND VPWR VPWR VGND _10129_/X hold512/A _10612_/S hold541/A sky130_fd_sc_hd__mux2_1
X_14937_ hold948/A _14937_/CLK _14937_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14868_ _14868_/Q _14868_/CLK _14868_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13787__904 VPWR VGND VPWR VGND _15159_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_07340_ _07340_/X _07166_/B _15472_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_14799_ _14799_/Q _14799_/CLK _14799_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09010_ VPWR VGND VGND VPWR _09890_/A _09010_/B _09010_/Y sky130_fd_sc_hd__nor2_1
X_07271_ VPWR VGND VGND VPWR _07272_/C _08041_/A _07271_/B sky130_fd_sc_hd__or2_1
XFILLER_31_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13828__945 VPWR VGND VPWR VGND _15200_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
Xhold157 hold157/X hold157/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/X hold168/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ VPWR VGND VGND VPWR _09931_/B _09917_/A _09912_/A sky130_fd_sc_hd__nor2_2
Xfanout615 VGND VPWR _11492_/S _11480_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout604 VPWR VGND _08411_/S _08409_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xhold179 hold179/X hold179/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout626 _09795_/S _09764_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout648 VPWR VGND _09552_/S _09521_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_09843_ VGND VPWR VPWR VGND _14179_/D hold480/X _09864_/S fanout61/X sky130_fd_sc_hd__mux2_1
Xfanout637 VPWR VGND _09617_/S _09591_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_13380__497 VPWR VGND VPWR VGND _14655_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_13988__1105 VPWR VGND VPWR VGND _15360_/CLK clkload19/A sky130_fd_sc_hd__inv_2
Xfanout659 VPWR VGND _09327_/S _09342_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09774_ VGND VPWR VPWR VGND _14275_/D fanout60/X _09795_/S hold507/X sky130_fd_sc_hd__mux2_1
X_08725_ VGND VPWR VGND VPWR _15271_/D hold976/X _08731_/A2 _08724_/X _11294_/A sky130_fd_sc_hd__o211a_1
X_08656_ VPWR VGND VGND VPWR _08655_/X _08690_/S _08194_/Y _14405_/Q _08656_/X _08654_/X
+ sky130_fd_sc_hd__o221a_1
X_08587_ VPWR VGND VPWR VGND _08586_/Y _10060_/C _08585_/Y _08992_/B _07534_/B sky130_fd_sc_hd__a22o_1
X_07607_ VPWR VGND VGND VPWR _07607_/C _07607_/B _07612_/A _07607_/Y sky130_fd_sc_hd__nor3_1
X_07538_ VPWR VGND VGND VPWR _07559_/A _07555_/A _07555_/B sky130_fd_sc_hd__or2_1
XFILLER_74_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13274__391 VPWR VGND VPWR VGND _14549_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_50_760 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_35_1327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07469_ VGND VPWR VPWR VGND _07471_/B _09311_/B _07469_/S _15593_/Q sky130_fd_sc_hd__mux2_1
XFILLER_22_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10480_ VPWR VGND VGND VPWR _10480_/X hold180/A _10484_/B sky130_fd_sc_hd__or2_1
X_09208_ VGND VPWR VPWR VGND _14885_/D hold1017/X _09213_/S clone55/A sky130_fd_sc_hd__mux2_1
XFILLER_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09139_ VGND VPWR VPWR VGND _14959_/D fanout62/X _09160_/S hold729/X sky130_fd_sc_hd__mux2_1
X_12150_ VPWR VGND VGND VPWR _12150_/X hold457/A _12155_/S sky130_fd_sc_hd__or2_1
X_11101_ VPWR VGND VPWR VGND _11098_/X _11112_/A _11100_/X _11101_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_300 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold680 hold680/X hold680/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13621__738 VPWR VGND VPWR VGND _14961_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_12081_ VGND VPWR VPWR VGND _12081_/X hold712/A _12227_/S hold238/A sky130_fd_sc_hd__mux2_1
XFILLER_78_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold691 hold691/X hold691/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ VGND VPWR VPWR VGND _11032_/X _11031_/X _11176_/S _11030_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1391 hold1391/X _15067_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1380 _09243_/A _14799_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14722_ hold454/A _14722_/CLK _14722_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11934_ VGND VPWR VGND VPWR _11934_/X _11931_/X _11933_/X _12156_/A1 _12212_/A1 sky130_fd_sc_hd__a211o_1
X_14653_ hold376/A _14653_/CLK _14653_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_587 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13515__632 VPWR VGND VPWR VGND _14790_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_60_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11865_ VPWR VGND VGND VPWR _11865_/X hold506/A _11882_/S sky130_fd_sc_hd__or2_1
X_11796_ VGND VPWR VPWR VGND _11796_/X _11793_/X _12591_/S _11792_/X sky130_fd_sc_hd__mux2_1
X_10816_ VPWR VGND VGND VPWR _10816_/X _10816_/A _10816_/B sky130_fd_sc_hd__or2_1
X_14584_ hold260/A _14584_/CLK _14584_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_484 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10747_ VPWR VGND VPWR VGND _10746_/X _10729_/A _11973_/B _10747_/X sky130_fd_sc_hd__a21o_1
X_10678_ VPWR VGND VGND VPWR _10678_/X hold231/A _10687_/B sky130_fd_sc_hd__or2_1
X_15205_ hold478/A _15205_/CLK _15205_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12417_ VPWR VGND VPWR VGND _12416_/X _12732_/A _12750_/B1 _12417_/X sky130_fd_sc_hd__a21o_1
X_12348_ VGND VPWR VGND VPWR _12348_/X _12345_/X _12347_/X _12375_/S _12376_/B2 sky130_fd_sc_hd__a211o_1
X_15136_ _15136_/Q _15136_/CLK _15136_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12279_ VGND VPWR VPWR VGND _12283_/B hold438/A _12689_/S hold268/A sky130_fd_sc_hd__mux2_1
X_15067_ _15067_/Q clkload14/A _15067_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_4_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_68_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_1314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08510_ VPWR VGND _15331_/D _08510_/B _08735_/C VPWR VGND sky130_fd_sc_hd__and2_1
X_09490_ VGND VPWR VPWR VGND _14569_/D fanout85/X _09514_/S hold415/X sky130_fd_sc_hd__mux2_1
XFILLER_3_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08441_ VGND VPWR VGND VPWR _15356_/D _15355_/Q _08448_/B _08440_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
X_13258__375 VPWR VGND VPWR VGND _14533_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_08372_ VGND VPWR VPWR VGND _15401_/D hold530/X _08372_/S _09228_/A0 sky130_fd_sc_hd__mux2_1
X_07323_ VPWR VGND VPWR VGND _07163_/A _07158_/Y _07159_/A _07323_/Y sky130_fd_sc_hd__a21oi_1
X_14034__1151 VPWR VGND VPWR VGND _15406_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_07254_ VPWR VGND VPWR VGND _07254_/Y _08066_/A sky130_fd_sc_hd__inv_2
XFILLER_69_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07185_ _07186_/B _15461_/Q _07345_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_2_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout401 VPWR VGND _11112_/A _10816_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout423 VPWR VGND _11104_/B1 fanout424/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout412 VGND VPWR _08178_/A1 _10717_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13963__1080 VPWR VGND VPWR VGND _15335_/CLK clkload28/A sky130_fd_sc_hd__inv_2
Xfanout456 VPWR VGND VGND VPWR clone2/A _10728_/S sky130_fd_sc_hd__buf_12
Xfanout445 VGND VPWR _11173_/A _11247_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1236 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout434 VPWR VGND _10930_/C1 _10891_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout489 VGND VPWR _11882_/S _12183_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09826_ VGND VPWR VPWR VGND _14226_/D _09826_/A1 _09833_/S hold213/X sky130_fd_sc_hd__mux2_1
Xfanout478 VGND VPWR _12089_/S _12097_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_12893__10 VPWR VGND VPWR VGND _14135_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_09757_ VGND VPWR VPWR VGND _14289_/D _09827_/A1 _09757_/S hold152/X sky130_fd_sc_hd__mux2_1
X_08708_ VGND VPWR VGND VPWR _08708_/X _14389_/Q _08664_/B _08711_/B1 _08654_/X sky130_fd_sc_hd__o211a_1
X_09688_ VGND VPWR VPWR VGND _14352_/D hold779/X _09693_/S _09688_/A0 sky130_fd_sc_hd__mux2_1
X_08639_ VGND VPWR VGND VPWR _08700_/A2 _14384_/Q _08194_/B _08639_/X sky130_fd_sc_hd__o21ba_1
X_11650_ VGND VPWR VPWR VGND _11654_/B hold666/A _11950_/B hold257/A sky130_fd_sc_hd__mux2_1
XFILLER_80_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_74_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout74 VPWR VGND VGND VPWR clone47/A fanout74/X sky130_fd_sc_hd__buf_8
Xfanout41 VPWR VGND fanout41/X clone6/A VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout63 VGND VPWR fanout63/X _07700_/X VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_11581_ VGND VPWR VGND VPWR _11581_/X _12099_/A1 _11577_/X _11580_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
Xfanout52 VPWR VGND VGND VPWR clone46/A fanout52/X sky130_fd_sc_hd__buf_8
X_10601_ VGND VPWR VPWR VGND _10605_/B hold521/A _10602_/S hold667/A sky130_fd_sc_hd__mux2_1
Xfanout85 VPWR VGND fanout85/X fanout86/X VPWR VGND sky130_fd_sc_hd__buf_6
X_10532_ VGND VPWR VPWR VGND _10532_/X hold735/A _10627_/S hold307/A sky130_fd_sc_hd__mux2_1
Xfanout96 VPWR VGND fanout96/X _08299_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_10463_ VGND VPWR VPWR VGND _10463_/X _14197_/Q _10464_/S hold478/A sky130_fd_sc_hd__mux2_1
X_13051__168 VPWR VGND VPWR VGND _14294_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_10394_ VPWR VGND VPWR VGND _10393_/X _10693_/B1 _10392_/X _10394_/Y sky130_fd_sc_hd__a21oi_1
X_12202_ VGND VPWR VGND VPWR _12202_/X _12230_/A1 _12198_/X _12201_/X _12202_/C1 sky130_fd_sc_hd__o211a_1
X_12133_ VGND VPWR VPWR VGND _12133_/X _14202_/Q _12155_/S hold328/A sky130_fd_sc_hd__mux2_1
XFILLER_46_1220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12064_ VPWR VGND VPWR VGND _12063_/X _12230_/C1 _12062_/X _12064_/Y sky130_fd_sc_hd__a21oi_1
X_11015_ VPWR VGND VPWR VGND _11014_/X _11023_/A1 _11013_/X _11015_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_58_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_61_800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14705_ hold491/A _14705_/CLK _14705_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_46_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11917_ VGND VPWR VPWR VGND _11918_/B _11916_/Y _12139_/S _11908_/Y sky130_fd_sc_hd__mux2_1
X_11848_ VPWR VGND VGND VPWR _11848_/X hold411/A _12089_/S sky130_fd_sc_hd__or2_1
X_14636_ hold460/A _14636_/CLK _14636_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14567_ hold456/A _14567_/CLK _14567_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13987__1104 VPWR VGND VPWR VGND _15359_/CLK clkload19/A sky130_fd_sc_hd__inv_2
X_11779_ VGND VPWR VPWR VGND _11779_/X hold473/A _12205_/S hold314/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1388 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14498_ hold787/A _14498_/CLK _14498_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_62_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkload22 VGND VPWR VGND VPWR clkload22/A clkload22/Y sky130_fd_sc_hd__bufinv_8
Xclkload44 clkload44/Y clkload44/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload33 clkload33/Y clkload33/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload11 clkload11/Y clkload11/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload55 VPWR VGND VPWR VGND clkload55/Y clkload55/A sky130_fd_sc_hd__inv_6
X_15119_ _15119_/Q _15119_/CLK _15119_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13643__760 VPWR VGND VPWR VGND _14983_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_08990_ VGND VPWR VGND VPWR _08990_/X _09873_/A _09016_/B1 _15106_/Q _08989_/Y sky130_fd_sc_hd__a211o_1
X_07941_ VPWR VGND VGND VPWR _07966_/A _07941_/Y _12813_/B sky130_fd_sc_hd__nand2_1
X_07872_ VPWR VGND VPWR VGND _15142_/Q clone18/X _07872_/Y _15353_/Q _08495_/A2 sky130_fd_sc_hd__a22oi_2
XFILLER_56_605 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09611_ VGND VPWR VPWR VGND _14457_/D _09625_/S fanout23/X hold1182/X sky130_fd_sc_hd__mux2_4
XFILLER_37_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09542_ VGND VPWR VPWR VGND _14520_/D fanout21/X _09553_/S hold155/X sky130_fd_sc_hd__mux2_1
X_09473_ VGND VPWR VPWR VGND _14583_/D fanout16/X _09485_/S hold307/X sky130_fd_sc_hd__mux2_1
X_08424_ VPWR VGND VGND VPWR _08425_/A _09937_/A _08424_/Y sky130_fd_sc_hd__nor2_1
X_08355_ VGND VPWR VPWR VGND _15418_/D hold786/X _08356_/S fanout45/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1357 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkload5 VGND VPWR VPWR VGND clkload5/A clkload5/Y sky130_fd_sc_hd__clkinvlp_4
X_07306_ VPWR VGND VGND VPWR _15465_/Q _07306_/B _07307_/B sky130_fd_sc_hd__nor2_1
X_08286_ VPWR VGND VGND VPWR _08286_/A _08286_/B _08286_/Y _10074_/S sky130_fd_sc_hd__nand3_1
X_07237_ VPWR VGND VPWR VGND _08199_/B _08201_/A _07213_/X _08179_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_1021 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07168_ VPWR VGND VGND VPWR _14405_/Q _07142_/X _07301_/B1 _07319_/B sky130_fd_sc_hd__o21a_1
X_07099_ VPWR VGND VPWR VGND _08290_/A _15445_/Q sky130_fd_sc_hd__inv_2
Xfanout231 VGND VPWR _12572_/C1 _12748_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout220 VGND VPWR fanout234/X _12115_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout253 VPWR VGND _12222_/C1 _07936_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout242 VGND VPWR _07955_/Y _08270_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout264 VGND VPWR _12029_/A _12103_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13692__809 VPWR VGND VPWR VGND _15032_/CLK clkload7/A sky130_fd_sc_hd__inv_2
Xfanout275 VGND VPWR fanout282/X _10583_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout297 VGND VPWR _10472_/S _10696_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout286 VGND VPWR _10604_/S _10612_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09809_ VGND VPWR VPWR VGND _14243_/D fanout60/X _09830_/S hold223/X sky130_fd_sc_hd__mux2_1
X_12820_ VPWR VGND VGND VPWR _12820_/A _12820_/Y _12820_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12751_ VPWR VGND VGND VPWR _12732_/Y _12750_/X _12751_/A2 _15476_/Q _15476_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
XFILLER_70_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12682_ VPWR VGND VGND VPWR _12682_/X _12698_/S _12682_/B sky130_fd_sc_hd__or2_1
X_15470_ _15470_/Q clkload38/A _15470_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11702_ VGND VPWR VPWR VGND _11702_/X _14865_/Q _12052_/S hold530/A sky130_fd_sc_hd__mux2_1
X_14421_ hold766/A _14421_/CLK _14421_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13586__703 VPWR VGND VPWR VGND _14917_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_11633_ VGND VPWR VPWR VGND _11633_/X _15482_/Q _12117_/B hold250/A sky130_fd_sc_hd__mux2_1
X_11564_ VPWR VGND VPWR VGND _11563_/Y _11280_/B _11542_/A _15442_/D sky130_fd_sc_hd__a21oi_1
XFILLER_10_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14352_ hold779/A _14352_/CLK _14352_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11495_ VGND VPWR VPWR VGND _15082_/D _11494_/X _11538_/S hold1405/X sky130_fd_sc_hd__mux2_1
X_14283_ hold563/A _14283_/CLK _14283_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10515_ VGND VPWR VGND VPWR _10515_/X _10634_/C1 _10510_/X _10514_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_13_1252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13627__744 VPWR VGND VPWR VGND _14967_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XFILLER_7_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10446_ VPWR VGND VGND VPWR _10446_/X _10557_/A _10446_/B sky130_fd_sc_hd__or2_1
X_10377_ VPWR VGND VPWR VGND _10376_/X _10618_/A _12121_/B1 _10377_/X sky130_fd_sc_hd__a21o_1
X_12116_ VGND VPWR VPWR VGND _12116_/X hold407/A _12117_/B hold736/A sky130_fd_sc_hd__mux2_1
X_12047_ VPWR VGND VPWR VGND _12046_/X _12103_/A _12047_/B1 _12047_/X sky130_fd_sc_hd__a21o_1
X_14033__1150 VPWR VGND VPWR VGND _15405_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
XFILLER_4_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14619_ hold639/A _14619_/CLK _14619_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15599_ VGND VPWR VGND VPWR _15599_/Q _15599_/D clkload55/A sky130_fd_sc_hd__dfxtp_4
X_08140_ VGND VPWR VGND VPWR _08140_/X _08182_/S _12774_/B _08139_/X _08280_/B2 sky130_fd_sc_hd__o211a_1
XFILLER_14_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_1152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_1065 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08071_ VGND VPWR VPWR VGND _15525_/D fanout17/X _08300_/S hold352/X sky130_fd_sc_hd__mux2_1
X_13073__190 VPWR VGND VPWR VGND _14316_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_08973_ VGND VPWR VGND VPWR _15113_/D hold791/X _08985_/A2 _08972_/X _08943_/A sky130_fd_sc_hd__o211a_1
X_07924_ VGND VPWR VGND VPWR _07924_/X _07984_/S _07918_/Y _07923_/Y _10071_/A sky130_fd_sc_hd__o211a_1
XFILLER_69_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13420__537 VPWR VGND VPWR VGND _14695_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_07855_ VPWR VGND VPWR VGND _07855_/B _07878_/B _07859_/A _07856_/B sky130_fd_sc_hd__or3_1
X_07786_ VPWR VGND VPWR VGND _08076_/B _07743_/B _07741_/X _08057_/A sky130_fd_sc_hd__a21o_1
XFILLER_37_660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09525_ VGND VPWR VPWR VGND _14537_/D fanout83/X _09537_/S hold210/X sky130_fd_sc_hd__mux2_1
XFILLER_40_803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk _12957__74/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09456_ VGND VPWR VPWR VGND _14600_/D clone49/A _09467_/S hold403/X sky130_fd_sc_hd__mux2_1
X_08407_ VGND VPWR VPWR VGND _15370_/D _09689_/A0 _08408_/S hold755/X sky130_fd_sc_hd__mux2_1
X_09387_ VGND VPWR VPWR VGND _14662_/D _09408_/S hold1128/X fanout74/X sky130_fd_sc_hd__mux2_4
X_13314__431 VPWR VGND VPWR VGND _14589_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_08338_ VGND VPWR VPWR VGND _15481_/D fanout96/X _08338_/S hold956/X sky130_fd_sc_hd__mux2_1
X_08269_ VPWR VGND VPWR VGND _08174_/Y _14836_/Q _08268_/X _08269_/Y sky130_fd_sc_hd__a21oi_1
X_11280_ VPWR VGND VPWR VGND _11567_/C _15443_/Q _11280_/B sky130_fd_sc_hd__or2_2
X_10300_ VGND VPWR VPWR VGND _10300_/X hold473/A _10664_/S hold314/A sky130_fd_sc_hd__mux2_1
X_10231_ VGND VPWR VPWR VGND _10235_/B hold746/A _10258_/B hold429/A sky130_fd_sc_hd__mux2_1
X_10162_ VGND VPWR VPWR VGND _10162_/X hold414/A _10484_/B hold200/A sky130_fd_sc_hd__mux2_1
X_14970_ hold406/A _14970_/CLK _14970_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10093_ VGND VPWR VPWR VGND _10093_/X _14187_/Q _10602_/S hold224/A sky130_fd_sc_hd__mux2_1
X_13986__1103 VPWR VGND VPWR VGND _15358_/CLK clkload19/A sky130_fd_sc_hd__inv_2
XFILLER_75_799 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12803_ VPWR VGND VPWR VGND _12878_/C _08542_/Y _12802_/X _15558_/D sky130_fd_sc_hd__a21oi_1
X_12734_ VGND VPWR VPWR VGND _12734_/X _14378_/Q _12736_/B _14730_/Q sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk _12979__96/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_10995_ VGND VPWR VPWR VGND _10995_/X _10994_/X _10995_/S _10993_/X sky130_fd_sc_hd__mux2_1
X_15522_ hold191/A _15522_/CLK _15522_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1038 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15453_ VGND VPWR VGND VPWR _15453_/Q _15453_/D clkload27/A sky130_fd_sc_hd__dfxtp_4
X_12665_ VGND VPWR VPWR VGND _12665_/X _12664_/X _12665_/S _12663_/X sky130_fd_sc_hd__mux2_1
X_12596_ VGND VPWR VGND VPWR _12596_/X _12593_/X _12595_/X _12748_/A1 _12596_/C1 sky130_fd_sc_hd__a211o_1
X_15384_ hold599/A _15384_/CLK _15384_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14404_ _14404_/Q clkload38/A _14404_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11616_ VGND VPWR VPWR VGND _11616_/X hold520/A _12097_/S hold309/A sky130_fd_sc_hd__mux2_1
X_13057__174 VPWR VGND VPWR VGND _14300_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_11547_ VGND VPWR _11545_/B hold1275/X _11547_/Y _15433_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
X_13942__1059 VPWR VGND VPWR VGND _15314_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_14335_ hold829/A _14335_/CLK _14335_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13861__978 VPWR VGND VPWR VGND _15233_/CLK clkload51/A sky130_fd_sc_hd__inv_2
Xhold509 hold509/X hold509/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ VGND VPWR VPWR VGND _11478_/X _15078_/Q _11490_/S _15076_/Q sky130_fd_sc_hd__mux2_1
X_14266_ hold645/A _14266_/CLK _14266_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14197_ _14197_/Q _14197_/CLK _14197_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10429_ VGND VPWR VGND VPWR _10429_/X hold730/A _10744_/A2 _10428_/X _10588_/S sky130_fd_sc_hd__o211a_1
XFILLER_48_1178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1209 hold1209/X _14130_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13755__872 VPWR VGND VPWR VGND _15127_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_07640_ VPWR VGND VGND VPWR _07640_/A _07972_/B _07640_/Y sky130_fd_sc_hd__nor2_1
X_07571_ VPWR VGND VGND VPWR _07573_/B _15445_/Q _07571_/B sky130_fd_sc_hd__or2_1
XFILLER_19_682 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clkload39/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09310_ VGND VPWR VPWR VGND _14731_/D fanout97/X _09310_/S hold165/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09241_ VPWR VGND VGND VPWR _09799_/B _09241_/Y _09694_/A sky130_fd_sc_hd__nor2_2
XFILLER_22_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09172_ VGND VPWR VPWR VGND _14919_/D hold386/X _09191_/S fanout64/X sky130_fd_sc_hd__mux2_1
X_08123_ _08128_/A _08120_/X _08121_/X _08122_/X _08294_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_30_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08054_ VGND VPWR VPWR VGND _08214_/B _08053_/X _08195_/A _07631_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08956_ VPWR VGND VGND VPWR _08983_/A _08956_/B _08956_/Y sky130_fd_sc_hd__nor2_1
X_08887_ VGND VPWR VGND VPWR _15149_/D hold1276/X _08893_/A2 _08886_/X _11974_/C1
+ sky130_fd_sc_hd__o211a_1
X_07907_ VGND VPWR VGND VPWR _07904_/X _07886_/A _12820_/A _07907_/X _07974_/B1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07838_ VPWR VGND _08023_/A _08022_/B _15557_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_72_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_clk clkload53/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07769_ VPWR VGND VGND VPWR _07769_/A _07769_/B _07770_/B _07769_/C sky130_fd_sc_hd__nand3_1
X_09508_ VGND VPWR VPWR VGND _14551_/D fanout16/X _09520_/S hold735/X sky130_fd_sc_hd__mux2_1
X_10780_ VGND VPWR VGND VPWR _10780_/X hold770/A _11215_/A2 _10779_/X _10315_/S sky130_fd_sc_hd__o211a_1
X_09439_ VGND VPWR VPWR VGND _14613_/D fanout8/X _09449_/S hold554/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12450_ VGND VPWR VGND VPWR _12450_/X _15504_/Q _12669_/A2 _12624_/S _12449_/X sky130_fd_sc_hd__o211a_1
X_11401_ VPWR VGND VPWR VGND _14852_/Q _14854_/Q _14853_/Q _11401_/Y _14851_/Q sky130_fd_sc_hd__nand4_1
X_12381_ VGND VPWR VGND VPWR _15466_/D _12491_/B1 _12379_/X _12380_/X _11567_/A sky130_fd_sc_hd__o211a_1
XANTENNA_91 _14385_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_80 fanout844/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_10_1200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11332_ VGND VPWR VPWR VGND _14830_/Q _11332_/X _14829_/Q sky130_fd_sc_hd__xor2_1
X_11263_ VGND VPWR VGND VPWR _11263_/X _11260_/X _11262_/X _10816_/A _11263_/C1 sky130_fd_sc_hd__a211o_1
X_13698__815 VPWR VGND VPWR VGND _15038_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_11194_ VGND VPWR VPWR VGND _11194_/X hold903/A _11204_/S hold594/A sky130_fd_sc_hd__mux2_1
X_10214_ VGND VPWR VPWR VGND _10214_/X _10213_/X _10995_/S _10212_/X sky130_fd_sc_hd__mux2_1
X_10145_ VGND VPWR VGND VPWR _10145_/X _10616_/A1 _10144_/X _10141_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
X_13739__856 VPWR VGND VPWR VGND _15111_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_14953_ hold808/A _14953_/CLK _14953_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_733 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10076_ VGND VPWR VGND VPWR _10075_/Y _10074_/X _15584_/Q _10072_/B _10075_/B _10076_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_78_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14884_ hold966/A _14884_/CLK _14884_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_758 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_clk clkload44/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_10978_ VPWR VGND VPWR VGND _10977_/X _11237_/A1 _10976_/X _10978_/Y sky130_fd_sc_hd__a21oi_1
X_12717_ VGND VPWR VPWR VGND _12717_/X _14346_/Q _12726_/S _15258_/Q sky130_fd_sc_hd__mux2_1
X_15505_ _15505_/Q _15505_/CLK _15505_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15436_ _15436_/Q clkload52/A _15436_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_31_666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12648_ VPWR VGND VPWR VGND _12647_/X _12656_/A1 _12646_/X _12648_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_699 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12579_ VPWR VGND VGND VPWR _12579_/X _12581_/S _12579_/B sky130_fd_sc_hd__or2_1
XFILLER_8_862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15367_ hold704/A _15367_/CLK _15367_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold317 hold317/X hold317/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold306 hold306/X hold306/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ _15298_/Q _15298_/CLK _15298_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14318_ hold476/A _14318_/CLK _14318_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14249_ hold377/A _14249_/CLK _14249_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold328 hold328/X hold328/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 hold339/X hold339/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout808 VPWR VGND _11399_/A1 _11398_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout819 VGND VPWR fanout824/X _11974_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_08810_ VGND VPWR VPWR VGND _15199_/D _09863_/A0 _08811_/S hold264/X sky130_fd_sc_hd__mux2_1
X_09790_ VGND VPWR VPWR VGND _14259_/D _09825_/A1 _09790_/S hold951/X sky130_fd_sc_hd__mux2_1
Xhold1006 hold1006/X _14491_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ VPWR VGND _15260_/D _08741_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
Xhold1017 hold1017/X _14885_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 hold1039/X _14499_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1028 hold1028/X _15494_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08672_ VGND VPWR VPWR VGND _08672_/X _14401_/Q _08684_/S _14385_/Q sky130_fd_sc_hd__mux2_1
XFILLER_6_1367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13491__608 VPWR VGND VPWR VGND _14766_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_07623_ VGND VPWR _07622_/X _07984_/S _07623_/Y _07621_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_18_clk clkload25/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07554_ VGND VPWR VGND VPWR _07555_/A _07560_/C _07554_/D _07558_/A _07555_/B sky130_fd_sc_hd__and4bb_4
X_07485_ VGND VPWR VGND VPWR _07486_/C _07580_/B _07580_/A _07577_/A _07483_/A sky130_fd_sc_hd__o211a_1
X_13532__649 VPWR VGND VPWR VGND _14863_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_09224_ VGND VPWR VPWR VGND _14869_/D hold827/X _09231_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_13985__1102 VPWR VGND VPWR VGND _15357_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_09155_ VGND VPWR VPWR VGND _14943_/D _09685_/A0 _09163_/S hold835/X sky130_fd_sc_hd__mux2_1
X_13385__502 VPWR VGND VPWR VGND _14660_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_14012__1129 VPWR VGND VPWR VGND _15384_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_09086_ VGND VPWR VPWR VGND _15007_/D hold1066/X _09094_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
X_08106_ VGND VPWR VGND VPWR _08106_/X _08280_/A2 _08103_/X _08102_/A _08105_/X sky130_fd_sc_hd__a211o_1
X_08037_ VGND VPWR _08037_/B _08037_/Y _08037_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13426__543 VPWR VGND VPWR VGND _14701_/CLK clkload23/A sky130_fd_sc_hd__inv_2
Xhold862 hold862/X hold862/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 hold840/X hold840/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 hold873/X hold873/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 hold851/X hold851/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 hold884/X hold884/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 hold895/X hold895/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09988_ VGND VPWR VPWR VGND _09988_/A _15610_/D _09989_/C sky130_fd_sc_hd__xor2_1
X_08939_ VPWR VGND _15128_/D _08939_/B _08955_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_44_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13941__1058 VPWR VGND VPWR VGND _15313_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_11950_ VPWR VGND VGND VPWR _11950_/X hold176/A _11950_/B sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_48_Left_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_714 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10901_ VPWR VGND VGND VPWR _10901_/X _11244_/S _10901_/B sky130_fd_sc_hd__or2_1
X_11881_ VGND VPWR VPWR VGND _11884_/B hold861/A _12183_/S hold710/A sky130_fd_sc_hd__mux2_1
X_10832_ VGND VPWR VPWR VGND _10832_/X hold573/A _11093_/S hold217/A sky130_fd_sc_hd__mux2_1
XFILLER_44_279 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10763_ VGND VPWR VPWR VGND _10763_/X _10760_/X _11092_/S _10759_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_482 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12502_ VGND VPWR VPWR VGND _12502_/X hold392/A _12539_/S hold370/A sky130_fd_sc_hd__mux2_1
X_12993__110 VPWR VGND VPWR VGND _14236_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_10694_ VPWR VGND VPWR VGND _10691_/X _10698_/A1 _10693_/X _10694_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_485 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15221_ hold285/A _15221_/CLK _15221_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_32_50 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12433_ VGND VPWR VPWR VGND _12433_/X _12430_/X _12536_/S _12429_/X sky130_fd_sc_hd__mux2_1
X_12364_ VGND VPWR VPWR VGND _12364_/X hold769/A _12370_/S hold475/A sky130_fd_sc_hd__mux2_1
X_15152_ _15152_/Q _15152_/CLK _15152_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11315_ VPWR VGND _14824_/D hold1292/X _11303_/A _11315_/A1 _11355_/S VGND VPWR sky130_fd_sc_hd__a31o_1
X_15083_ _15083_/Q clkload37/A _15083_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_4_331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12295_ VGND VPWR VGND VPWR _12295_/X _12294_/X _12293_/X _12698_/S _12702_/C1 sky130_fd_sc_hd__a211o_1
X_13169__286 VPWR VGND VPWR VGND _14444_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_11246_ VGND VPWR VPWR VGND _11247_/B _11245_/Y _11246_/S _11237_/Y sky130_fd_sc_hd__mux2_1
X_11177_ VPWR VGND VGND VPWR _11177_/X hold424/A _11179_/S sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_66_Left_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10128_ VGND VPWR VPWR VGND _10132_/B hold427/A _10612_/S hold548/A sky130_fd_sc_hd__mux2_1
X_10059_ VPWR VGND VGND VPWR _10059_/A _12878_/C _15640_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14936_ hold873/A _14936_/CLK _14936_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14867_ hold778/A _14867_/CLK _14867_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14798_ hold489/A _14798_/CLK _14798_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07270_ VPWR VGND VGND VPWR _08026_/A _08010_/A _08047_/A _07270_/Y sky130_fd_sc_hd__nor3_1
X_13867__984 VPWR VGND VPWR VGND _15239_/CLK clkload9/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_75_Left_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12969__86 VPWR VGND VPWR VGND _14212_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_15419_ hold475/A _15419_/CLK _15419_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13113__230 VPWR VGND VPWR VGND _14356_/CLK clkload17/A sky130_fd_sc_hd__inv_2
Xhold147 hold147/X hold147/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ VGND VPWR VGND VPWR _14140_/D _09931_/B _14140_/Q _09910_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_7_clk clkload13/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold158 hold158/X hold158/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 hold169/X hold169/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout605 VGND VPWR _08377_/Y _08409_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout638 _09619_/S _09622_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout616 VGND VPWR _11441_/Y _11492_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout627 _09763_/S _09756_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout649 VPWR VGND _09520_/S _09513_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09842_ VGND VPWR VPWR VGND _14180_/D hold642/X _09861_/S fanout65/X sky130_fd_sc_hd__mux2_1
XFILLER_8_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09773_ VGND VPWR VPWR VGND _14276_/D fanout66/X _09792_/S hold392/X sky130_fd_sc_hd__mux2_1
X_08724_ VPWR VGND VPWR VGND hold1451/X _08523_/B _08724_/X _08728_/B1 _14382_/Q _08726_/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_54_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08655_ VPWR VGND VGND VPWR _08655_/X _14389_/Q _08664_/B sky130_fd_sc_hd__or2_1
XFILLER_74_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08586_ VGND VPWR _08586_/B _08586_/Y _08586_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_53_27 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_42_706 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07606_ VGND VPWR VPWR VGND _07612_/A _07606_/X _07606_/B sky130_fd_sc_hd__xor2_1
X_07537_ VGND VPWR VGND VPWR _07555_/B _07552_/B1 _07533_/X _15566_/Q _07536_/X sky130_fd_sc_hd__a211o_1
XFILLER_35_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07468_ VPWR VGND VGND VPWR _07487_/A _07486_/A _07468_/B sky130_fd_sc_hd__nand2_1
X_07399_ _07665_/B _07397_/A _07397_/B _07397_/C _07398_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09207_ VGND VPWR VPWR VGND _14886_/D hold964/X _09228_/S fanout62/X sky130_fd_sc_hd__mux2_1
X_09138_ VGND VPWR VPWR VGND _14960_/D fanout64/X _09157_/S hold845/X sky130_fd_sc_hd__mux2_1
X_11100_ VPWR VGND VPWR VGND _11099_/X _11110_/A _11263_/C1 _11100_/X sky130_fd_sc_hd__a21o_1
X_09069_ VGND VPWR VPWR VGND _15024_/D hold1110/X _09090_/S fanout64/X sky130_fd_sc_hd__mux2_1
XFILLER_11_1372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold681 hold681/X hold681/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13660__777 VPWR VGND VPWR VGND _15000_/CLK clkload8/A sky130_fd_sc_hd__inv_2
Xhold670 hold670/X hold670/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12080_ VGND VPWR VGND VPWR _12080_/X _15494_/Q _12080_/A2 _12069_/S _12079_/X sky130_fd_sc_hd__o211a_1
X_11031_ VGND VPWR VPWR VGND _11031_/X hold955/A _11175_/S hold561/A sky130_fd_sc_hd__mux2_1
Xhold692 hold692/X hold692/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1370 hold1370/X _15062_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1392 hold1392/X _15323_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1381 _10002_/A _15616_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14721_ hold465/A _14721_/CLK _14721_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11933_ VGND VPWR VGND VPWR _11933_/X _15008_/Q _12229_/A2 _11925_/S _11932_/X sky130_fd_sc_hd__o211a_1
XFILLER_60_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11864_ VGND VPWR VPWR VGND _11864_/X hold806/A _11876_/B hold443/A sky130_fd_sc_hd__mux2_1
X_14652_ hold319/A _14652_/CLK _14652_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13554__671 VPWR VGND VPWR VGND _14885_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_10815_ VGND VPWR VGND VPWR _10815_/X _10816_/A _10811_/X _10814_/X _11259_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_45_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11795_ VGND VPWR VGND VPWR _11795_/X _12588_/A1 _11791_/X _11794_/X _12572_/C1 sky130_fd_sc_hd__o211a_1
X_14583_ hold307/A _14583_/CLK _14583_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10746_ VPWR VGND _10746_/X _10745_/X _10741_/X clone2/X _10737_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10677_ VGND VPWR VPWR VGND _10677_/X _10676_/X _10677_/S _10675_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_16_1283 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15204_ hold303/A _15204_/CLK _15204_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12416_ VPWR VGND _12416_/X _12415_/X _12411_/X _12731_/S _12407_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15135_ _15135_/Q _15135_/CLK _15135_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12347_ VGND VPWR VGND VPWR _12347_/X _14496_/Q _12861_/A1 _12367_/S _12346_/X sky130_fd_sc_hd__o211a_1
X_12278_ VPWR VGND VPWR VGND _12277_/X _12703_/A1 _12276_/X _12278_/Y sky130_fd_sc_hd__a21oi_1
X_15066_ _15066_/Q clkload14/A _15066_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11229_ VPWR VGND VGND VPWR _11210_/Y _11228_/X _12677_/A2 _14409_/Q _14409_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
X_13984__1101 VPWR VGND VPWR VGND _15356_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_3_1326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14919_ hold386/A _14919_/CLK _14919_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14011__1128 VPWR VGND VPWR VGND _15383_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_08440_ VPWR VGND VGND VPWR _08440_/X _15356_/Q _08488_/B sky130_fd_sc_hd__or2_1
X_08371_ VGND VPWR VPWR VGND _15402_/D hold556/X _08372_/S _09863_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_17_1003 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07322_ VGND VPWR VGND VPWR _07639_/A _07320_/X _07170_/Y _07663_/A _07663_/B _07619_/B
+ sky130_fd_sc_hd__a311o_1
X_07253_ VPWR VGND VPWR VGND _08066_/A _08041_/A _08067_/A sky130_fd_sc_hd__or2_2
X_13940__1057 VPWR VGND VPWR VGND _15312_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_07184_ VGND VPWR VGND VPWR _07186_/A _14395_/Q _07304_/A2 _07304_/B1 _15461_/Q sky130_fd_sc_hd__o211a_1
XFILLER_69_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout402 VGND VPWR _10846_/A1 _10816_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout413 VPWR VGND _10741_/C1 _08178_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout446 VPWR VGND _11173_/A _11210_/A VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout435 VGND VPWR _11023_/A1 _10891_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout424 VPWR VGND fanout424/X _07852_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout457 VPWR VGND _10987_/S clone2/A VPWR VGND sky130_fd_sc_hd__buf_4
X_09825_ VGND VPWR VPWR VGND _14227_/D _09825_/A1 _09825_/S hold197/X sky130_fd_sc_hd__mux2_1
X_13497__614 VPWR VGND VPWR VGND _14772_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
Xfanout479 VGND VPWR _12089_/S _11838_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout468 VGND VPWR _12861_/A1 _12488_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09756_ VGND VPWR VPWR VGND _14290_/D _09826_/A1 _09756_/S hold431/X sky130_fd_sc_hd__mux2_1
X_09687_ VGND VPWR VPWR VGND _14353_/D hold859/X _09687_/S _09792_/A1 sky130_fd_sc_hd__mux2_1
XFILLER_41_1387 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13538__655 VPWR VGND VPWR VGND _14869_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_08707_ VGND VPWR VGND VPWR _15279_/D hold1116/X _08721_/A2 _08706_/X _12159_/C1
+ sky130_fd_sc_hd__o211a_1
X_08638_ VGND VPWR VGND VPWR _15298_/D hold1007/X _08701_/A2 _08637_/X _12233_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_547 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08569_ VGND VPWR VGND VPWR _08569_/X _08605_/A _08615_/B1 hold1080/X _08568_/Y sky130_fd_sc_hd__a211o_1
Xfanout31 VPWR VGND fanout31/X fanout34/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout20 VGND VPWR _08051_/X fanout20/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout42 VPWR VGND VGND VPWR clone44/A fanout42/X sky130_fd_sc_hd__buf_8
Xfanout64 VPWR VGND fanout64/X fanout67/X VPWR VGND sky130_fd_sc_hd__buf_2
X_11580_ VPWR VGND VGND VPWR _11580_/X _12098_/A _11580_/B sky130_fd_sc_hd__or2_1
Xfanout53 VPWR VGND VGND VPWR clone5/A clone46/A sky130_fd_sc_hd__buf_8
X_10600_ VPWR VGND VGND VPWR _10581_/Y _10599_/X _10562_/B _14392_/Q _14392_/D _12085_/C1
+ sky130_fd_sc_hd__o221a_1
Xfanout75 VPWR VGND VGND VPWR _07659_/X clone47/A sky130_fd_sc_hd__buf_8
Xfanout86 VPWR VGND VGND VPWR _07614_/X fanout86/X sky130_fd_sc_hd__buf_8
X_10531_ VGND VPWR VGND VPWR _10531_/X hold850/A _10629_/A2 _10530_/X _10634_/A1 sky130_fd_sc_hd__o211a_1
Xfanout97 VPWR VGND fanout97/X _08299_/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_13_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xwire858 VGND VPWR wire858/X wire858/A VPWR VGND sky130_fd_sc_hd__buf_1
X_10462_ VGND VPWR VPWR VGND _10462_/X hold901/A _10464_/S hold176/A sky130_fd_sc_hd__mux2_1
X_12201_ VPWR VGND VGND VPWR _12201_/X _12221_/S _12201_/B sky130_fd_sc_hd__or2_1
X_10393_ VGND VPWR VPWR VGND _10393_/X _10390_/X _10685_/S _10389_/X sky130_fd_sc_hd__mux2_1
X_12132_ VGND VPWR VPWR VGND _12132_/X hold645/A _12155_/S hold621/A sky130_fd_sc_hd__mux2_1
X_12063_ VGND VPWR VPWR VGND _12063_/X _12060_/X _12221_/S _12059_/X sky130_fd_sc_hd__mux2_1
X_11014_ VGND VPWR VPWR VGND _11014_/X _11011_/X _11162_/S _11010_/X sky130_fd_sc_hd__mux2_1
X_14211__929 _14211_/D _14211__929/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_65_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14704_ hold494/A _14704_/CLK _14704_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11916_ VPWR VGND VPWR VGND _11915_/X _12230_/C1 _11914_/X _11916_/Y sky130_fd_sc_hd__a21oi_1
X_13290__407 VPWR VGND VPWR VGND _14565_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_11847_ VGND VPWR VPWR VGND _11847_/X _11846_/X _12100_/S _11845_/X sky130_fd_sc_hd__mux2_1
X_14635_ hold692/A _14635_/CLK _14635_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14566_ _14566_/Q _14566_/CLK _14566_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11778_ VGND VPWR VGND VPWR _11778_/X _12008_/C1 _11773_/X _11777_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_18_1334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_53_1258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13331__448 VPWR VGND VPWR VGND _14606_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_10729_ VPWR VGND VGND VPWR _10729_/A _10729_/B _10729_/Y sky130_fd_sc_hd__nor2_1
X_12939__56 VPWR VGND VPWR VGND _14182_/CLK clkload52/A sky130_fd_sc_hd__inv_2
X_14497_ _14497_/Q _14497_/CLK _14497_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkload23 clkload23/Y clkload23/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload12 VGND VPWR VGND VPWR clkload12/Y clkload12/A sky130_fd_sc_hd__inv_12
Xclkload34 VGND VPWR VPWR VGND clkload34/A clkload34/Y sky130_fd_sc_hd__clkinv_2
Xclkload45 VPWR VGND VGND VPWR clkload45/Y clkload45/A sky130_fd_sc_hd__inv_16
XFILLER_55_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15118_ hold988/A _15118_/CLK _15118_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13184__301 VPWR VGND VPWR VGND _14459_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_5_470 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15049_ hold432/A _15049_/CLK _15049_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07940_ VGND VPWR VPWR VGND _07945_/A _12813_/B _07940_/B sky130_fd_sc_hd__xor2_1
XFILLER_64_1354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13225__342 VPWR VGND VPWR VGND _14500_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_07871_ VGND VPWR VPWR VGND _15535_/D fanout54/X _08231_/S hold288/X sky130_fd_sc_hd__mux2_1
XFILLER_68_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09610_ VGND VPWR VPWR VGND _14458_/D fanout27/X _09617_/S hold566/X sky130_fd_sc_hd__mux2_1
XFILLER_7_1270 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_37_853 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09541_ VGND VPWR VPWR VGND _14521_/D fanout25/X _09555_/S hold202/X sky130_fd_sc_hd__mux2_1
XFILLER_37_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09472_ VGND VPWR VPWR VGND _14584_/D fanout20/X _09478_/S hold260/X sky130_fd_sc_hd__mux2_1
X_08423_ VPWR VGND VGND VPWR _14767_/Q _09937_/A _15365_/Q sky130_fd_sc_hd__nand2_1
X_08354_ VGND VPWR VPWR VGND _15419_/D hold475/X _08372_/S fanout50/X sky130_fd_sc_hd__mux2_1
X_07305_ VPWR VGND _07311_/B _07306_/B _15465_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_08285_ VGND VPWR VPWR VGND _15514_/D _09692_/A0 _08300_/S hold233/X sky130_fd_sc_hd__mux2_1
Xclkload6 VGND VPWR VPWR VGND clkload6/A clkload6/Y sky130_fd_sc_hd__clkinv_2
X_07236_ VPWR VGND VPWR VGND _08222_/B _08223_/A _07216_/X _08199_/B sky130_fd_sc_hd__a21o_1
X_07167_ VPWR VGND VPWR VGND _07167_/Y _07338_/B sky130_fd_sc_hd__inv_2
X_07098_ VPWR VGND VPWR VGND _07360_/A _15446_/Q sky130_fd_sc_hd__inv_2
X_12953__70 VPWR VGND VPWR VGND _14196_/CLK clkload18/A sky130_fd_sc_hd__inv_2
Xfanout221 VGND VPWR _12189_/C1 _12184_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout232 VGND VPWR _12572_/C1 _12702_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout210 VGND VPWR _12674_/A1 _12662_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout254 VPWR VGND _12740_/C1 _12864_/A1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout265 VPWR VGND _12029_/A _12214_/A VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout243 VPWR VGND _12722_/A1 _12376_/B2 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout298 VGND VPWR _10484_/B _10464_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout287 VGND VPWR _10604_/S _10353_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09808_ VGND VPWR VPWR VGND _14244_/D fanout65/X _09827_/S hold364/X sky130_fd_sc_hd__mux2_1
Xfanout276 VGND VPWR _12866_/A1 _11003_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09739_ VGND VPWR VPWR VGND _14307_/D fanout60/X _09760_/S hold293/X sky130_fd_sc_hd__mux2_1
X_13772__889 VPWR VGND VPWR VGND _15144_/CLK clkload23/A sky130_fd_sc_hd__inv_2
X_12750_ VPWR VGND VPWR VGND _12749_/X _12732_/A _12750_/B1 _12750_/X sky130_fd_sc_hd__a21o_1
X_12681_ VGND VPWR VPWR VGND _12681_/X hold415/A _12689_/S hold234/A sky130_fd_sc_hd__mux2_1
X_11701_ VGND VPWR VGND VPWR _11701_/X hold967/A _12488_/A2 _12489_/A1 _11700_/X sky130_fd_sc_hd__o211a_1
X_14420_ hold885/A _14420_/CLK _14420_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11632_ VGND VPWR VGND VPWR _11632_/X hold704/A _12040_/A2 _12008_/A1 _11631_/X sky130_fd_sc_hd__o211a_1
X_14351_ _14351_/Q _14351_/CLK _14351_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11563_ VPWR VGND VGND VPWR _11563_/A _11563_/Y _11563_/B sky130_fd_sc_hd__nand2_1
X_13666__783 VPWR VGND VPWR VGND _15006_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_11494_ VGND VPWR VPWR VGND _11494_/X _11493_/X _11537_/S _15462_/Q sky130_fd_sc_hd__mux2_1
X_14282_ _14282_/Q _14282_/CLK _14282_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10514_ VGND VPWR VGND VPWR _10514_/X _10513_/X _10512_/X _10510_/S _10630_/C1 sky130_fd_sc_hd__a211o_1
X_13983__1100 VPWR VGND VPWR VGND _15355_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_40_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10445_ VGND VPWR VGND VPWR _10445_/X _10557_/A _10441_/X _10444_/X _10717_/C1 sky130_fd_sc_hd__o211a_1
X_14010__1127 VPWR VGND VPWR VGND _15382_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_10376_ VPWR VGND _10376_/X _10375_/X _10371_/X _10617_/S _10367_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12115_ VGND VPWR VGND VPWR _12115_/X _12112_/X _12114_/X _12119_/A1 _12115_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_2_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13209__326 VPWR VGND VPWR VGND _14484_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_12046_ VPWR VGND _12046_/X _12045_/X _12041_/X _12176_/S _12037_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_77_296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_59_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_653 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12879_ VPWR VGND VPWR VGND _08194_/Y _07574_/A _12878_/X _15602_/D sky130_fd_sc_hd__a21oi_1
XFILLER_60_152 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14618_ hold515/A _14618_/CLK _14618_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15598_ VGND VPWR VGND VPWR _15598_/Q _15598_/D clkload45/A sky130_fd_sc_hd__dfxtp_4
X_14549_ hold877/A _14549_/CLK _14549_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08070_ VGND VPWR VPWR VGND _08070_/D _08070_/C _08070_/B _08070_/A _08070_/X sky130_fd_sc_hd__or4_4
X_14192__910 _14192_/D _14192__910/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08972_ VPWR VGND VGND VPWR _08972_/X _08972_/A _08972_/B sky130_fd_sc_hd__or2_1
X_07923_ VPWR VGND VGND VPWR _07984_/S _07923_/Y _07923_/B sky130_fd_sc_hd__nand2_1
X_07854_ VGND VPWR _07854_/B _12831_/B _07859_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07785_ VPWR VGND VPWR VGND _08097_/A _07745_/X _08096_/B _08076_/B sky130_fd_sc_hd__a21o_1
XFILLER_25_801 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09524_ _14538_/D fanout93/X fanout89/X _09522_/Y _09523_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_13002__119 VPWR VGND VPWR VGND _14245_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_09455_ VGND VPWR VPWR VGND _14601_/D fanout85/X _09467_/S hold234/X sky130_fd_sc_hd__mux2_1
X_08406_ VGND VPWR VPWR VGND _15371_/D _09550_/A1 _08411_/S hold473/X sky130_fd_sc_hd__mux2_1
X_13353__470 VPWR VGND VPWR VGND _14628_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_09386_ VGND VPWR VPWR VGND _14663_/D hold388/X _09408_/S fanout78/X sky130_fd_sc_hd__mux2_1
X_08337_ VGND VPWR VPWR VGND _15482_/D _09658_/A0 _08338_/S hold1002/X sky130_fd_sc_hd__mux2_1
X_08268_ VPWR VGND VPWR VGND clone20/X _15333_/Q _07567_/B _08268_/X _15154_/Q sky130_fd_sc_hd__a22o_1
X_07219_ VPWR VGND _07219_/X _07234_/B _15448_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_08199_ VGND VPWR _08199_/B _08200_/B _08201_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_10230_ VPWR VGND VGND VPWR _10211_/Y _10229_/X _12380_/B _14382_/Q _14382_/D _12085_/C1
+ sky130_fd_sc_hd__o221a_1
X_10161_ VGND VPWR VGND VPWR _10161_/X hold957/A _10688_/A2 _10160_/X _10486_/A1 sky130_fd_sc_hd__o211a_1
X_13700__817 VPWR VGND VPWR VGND _15040_/CLK clkload13/A sky130_fd_sc_hd__inv_2
XFILLER_10_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10092_ VGND VPWR VPWR VGND _10092_/X hold366/A _10602_/S hold563/A sky130_fd_sc_hd__mux2_1
XFILLER_78_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12802_ VPWR VGND VGND VPWR _10079_/X _08000_/Y _12820_/B _07999_/X _12802_/X _12801_/X
+ sky130_fd_sc_hd__o221a_1
X_10994_ VGND VPWR VPWR VGND _10994_/X hold776/A _10994_/S hold446/A sky130_fd_sc_hd__mux2_1
X_15521_ hold271/A _15521_/CLK _15521_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12733_ VGND VPWR VPWR VGND _12733_/X _14442_/Q _12736_/B _14698_/Q sky130_fd_sc_hd__mux2_1
XFILLER_43_686 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15452_ VGND VPWR VGND VPWR _15452_/Q _15452_/D clkload9/A sky130_fd_sc_hd__dfxtp_4
X_12664_ VGND VPWR VPWR VGND _12664_/X _14376_/Q _12664_/S _14728_/Q sky130_fd_sc_hd__mux2_1
X_14403_ _14403_/Q clkload36/A _14403_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12595_ VGND VPWR VGND VPWR _12595_/X _15026_/Q _12746_/A2 _12591_/S _12594_/X sky130_fd_sc_hd__o211a_1
X_11615_ VGND VPWR VPWR VGND _11615_/X _14188_/Q _12097_/S hold186/A sky130_fd_sc_hd__mux2_1
X_15383_ hold633/A _15383_/CLK _15383_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11546_ VPWR VGND VPWR VGND _11545_/Y _11271_/B _11542_/A _15433_/D sky130_fd_sc_hd__a21oi_1
X_14334_ _14334_/Q _14334_/CLK _14334_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12909__26 VPWR VGND VPWR VGND _14151_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_14265_ _14265_/Q _14265_/CLK _14265_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11477_ VGND VPWR VPWR VGND _15076_/D _11476_/X _11477_/S _15076_/Q sky130_fd_sc_hd__mux2_1
X_14217__935 _14217_/D _14217__935/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_14196_ _14196_/Q _14196_/CLK _14196_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10428_ VPWR VGND VGND VPWR _10428_/X hold292/A _10742_/S sky130_fd_sc_hd__or2_1
X_10359_ VPWR VGND VGND VPWR _10618_/A _10359_/B _10359_/Y sky130_fd_sc_hd__nor2_1
X_12029_ VPWR VGND VGND VPWR _12029_/A _12029_/B _12029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13296__413 VPWR VGND VPWR VGND _14571_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_07570_ VGND VPWR VPWR VGND _07570_/X _12080_/A2 _08195_/A _07561_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09240_ VPWR VGND VPWR VGND _09556_/C _09799_/B _09240_/A _09311_/B sky130_fd_sc_hd__or3b_2
X_13337__454 VPWR VGND VPWR VGND _14612_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_14125__1242 VPWR VGND VPWR VGND _15544_/CLK clkload54/A sky130_fd_sc_hd__inv_2
XFILLER_72_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09171_ VGND VPWR VPWR VGND _14920_/D hold764/X _09191_/S fanout68/X sky130_fd_sc_hd__mux2_1
X_08122_ VPWR VGND VPWR VGND _08278_/B _08116_/A _08280_/A2 _08122_/X _07244_/A sky130_fd_sc_hd__a22o_1
X_08053_ VPWR VGND VPWR VGND _08252_/A2 _15344_/Q _08253_/A2 _08053_/X _15149_/Q sky130_fd_sc_hd__a22o_1
X_12923__40 VPWR VGND VPWR VGND _14166_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_08955_ VPWR VGND _15119_/D _08955_/B _08955_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07906_ VPWR VGND VGND VPWR _12820_/A _07906_/A _07906_/B sky130_fd_sc_hd__or2_1
X_08886_ VPWR VGND VGND VPWR _08886_/X _15149_/Q _08918_/B sky130_fd_sc_hd__or2_1
X_07837_ VPWR VGND VPWR VGND _07837_/Y _08022_/B sky130_fd_sc_hd__inv_2
X_07768_ VPWR VGND VGND VPWR _14153_/Q _08273_/A _08272_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09507_ VGND VPWR VPWR VGND _14552_/D fanout20/X _09513_/S hold640/X sky130_fd_sc_hd__mux2_1
X_07699_ VPWR VGND VPWR VGND _07698_/X _15630_/Q _07929_/A2 _07699_/X _08249_/B2 sky130_fd_sc_hd__a22o_1
XFILLER_24_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09438_ VGND VPWR VPWR VGND _14614_/D fanout13/X _09449_/S hold916/X sky130_fd_sc_hd__mux2_1
X_09369_ VGND VPWR VPWR VGND _14677_/D hold849/X _09379_/S fanout10/X sky130_fd_sc_hd__mux2_1
XFILLER_36_1050 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11400_ VGND VPWR _11400_/B _14853_/D _11400_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_12380_ VPWR VGND VGND VPWR _12380_/X _15466_/Q _12380_/B sky130_fd_sc_hd__or2_1
X_11331_ VGND VPWR VGND VPWR _11330_/X _14829_/Q _11316_/Y _14829_/D sky130_fd_sc_hd__o21ba_1
XANTENNA_70 _09864_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_81 _07994_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_92 _14400_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_13130__247 VPWR VGND VPWR VGND _14373_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_11262_ VGND VPWR VGND VPWR _11262_/X _15030_/Q _11262_/A2 _11261_/X _10851_/A sky130_fd_sc_hd__o211a_1
XFILLER_21_74 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11193_ VGND VPWR VPWR VGND _11197_/B hold500/A _11216_/S hold577/A sky130_fd_sc_hd__mux2_1
X_10213_ VGND VPWR VPWR VGND _10213_/X _14350_/Q _10567_/S hold468/A sky130_fd_sc_hd__mux2_1
X_10144_ VGND VPWR VPWR VGND _10144_/X _10143_/X _10144_/S _10142_/X sky130_fd_sc_hd__mux2_1
X_13778__895 VPWR VGND VPWR VGND _15150_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_10075_ VPWR VGND VGND VPWR _10075_/A _10075_/B _10075_/Y sky130_fd_sc_hd__nor2_1
X_14952_ hold792/A _14952_/CLK _14952_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14883_ hold769/A _14883_/CLK _14883_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_918 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13024__141 VPWR VGND VPWR VGND _14267_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_1_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10977_ VGND VPWR VPWR VGND _10977_/X _10974_/X _10995_/S _10973_/X sky130_fd_sc_hd__mux2_1
X_12716_ VGND VPWR VPWR VGND _12716_/X _14506_/Q _12716_/S _14186_/Q sky130_fd_sc_hd__mux2_1
X_15504_ _15504_/Q _15504_/CLK _15504_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_16_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15435_ _15435_/Q clkload47/A _15435_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12647_ VGND VPWR VPWR VGND _12647_/X _12644_/X _12655_/S _12643_/X sky130_fd_sc_hd__mux2_1
X_15366_ hold931/A _15366_/CLK _15366_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12578_ VGND VPWR VPWR VGND _12578_/X _14470_/Q _12578_/S _14758_/Q sky130_fd_sc_hd__mux2_1
X_14317_ hold957/A _14317_/CLK _14317_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold307 hold307/X hold307/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11529_ VGND VPWR VPWR VGND _11529_/X _15095_/Q _11529_/S _15093_/Q sky130_fd_sc_hd__mux2_1
X_15297_ _15297_/Q _15297_/CLK _15297_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold329 hold329/X hold329/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 hold318/X hold318/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ hold276/A _14248_/CLK _14248_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14179_ hold480/A _14179_/CLK _14179_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout809 VGND VPWR _08529_/A _11398_/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_08740_ VPWR VGND VPWR VGND _09938_/C _14766_/Q _08522_/B _08741_/B _15260_/Q sky130_fd_sc_hd__a22o_1
Xhold1007 hold1007/X _15298_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 hold1018/X _14553_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 hold1029/X _14351_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08671_ VGND VPWR VGND VPWR _15291_/D hold1375/X _08701_/A2 _08670_/X _12085_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_1149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_597 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07622_ VPWR VGND VGND VPWR _07621_/B _07637_/A _07625_/A _07622_/X sky130_fd_sc_hd__o21a_1
X_07553_ VPWR VGND VGND VPWR _07560_/B _07560_/D _07554_/D sky130_fd_sc_hd__nor2_1
X_13571__688 VPWR VGND VPWR VGND _14902_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_07484_ VPWR VGND VGND VPWR _07580_/A _07580_/B _07483_/A _07578_/A sky130_fd_sc_hd__o21a_1
XFILLER_50_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_34_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09223_ VGND VPWR VPWR VGND _14870_/D hold910/X _09231_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_21_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09154_ VGND VPWR VPWR VGND _14944_/D fanout7/X _09161_/S hold525/X sky130_fd_sc_hd__mux2_1
X_08105_ VPWR VGND VPWR VGND _15075_/Q _11440_/B _08105_/X _08293_/A3 _07195_/A _08104_/Y
+ sky130_fd_sc_hd__a221o_1
X_09085_ VGND VPWR VPWR VGND _15008_/D hold1024/X _09092_/S fanout5/X sky130_fd_sc_hd__mux2_1
Xhold830 hold830/X hold830/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08036_ VPWR VGND VGND VPWR _08035_/X _07421_/Y _08034_/X _07421_/A _08051_/A _07996_/X
+ sky130_fd_sc_hd__o221a_1
Xhold852 hold852/X hold852/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 hold841/X hold841/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold863 hold863/X hold863/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13465__582 VPWR VGND VPWR VGND _14740_/CLK clkload18/A sky130_fd_sc_hd__inv_2
Xhold896 hold896/X hold896/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 hold874/X hold874/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 hold885/X hold885/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09987_ VPWR VGND VGND VPWR _09989_/C _09987_/B _15609_/D sky130_fd_sc_hd__nor2_1
X_08938_ VPWR VGND VPWR VGND _08969_/A _15127_/Q _08933_/A _08938_/X hold1412/X sky130_fd_sc_hd__a22o_1
XFILLER_40_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13008__125 VPWR VGND VPWR VGND _14251_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_08869_ VGND VPWR VGND VPWR _08869_/X hold1253/X _08893_/A2 _08868_/X _09024_/A sky130_fd_sc_hd__o211a_1
XFILLER_79_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_214 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10900_ VGND VPWR VPWR VGND _10900_/X _14561_/Q _10919_/S _14593_/Q sky130_fd_sc_hd__mux2_1
X_13812__929 VPWR VGND VPWR VGND _15184_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_11880_ VGND VPWR VPWR VGND _11880_/X hold933/A _12183_/S hold686/A sky130_fd_sc_hd__mux2_1
X_10831_ VGND VPWR VPWR VGND _10831_/X _14207_/Q _11093_/S hold274/A sky130_fd_sc_hd__mux2_1
X_10762_ VGND VPWR VGND VPWR _10762_/X _11086_/C1 _10758_/X _10761_/X _11104_/B1 sky130_fd_sc_hd__o211a_1
XFILLER_25_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12501_ VGND VPWR VPWR VGND _12505_/B hold560/A _12539_/S hold364/A sky130_fd_sc_hd__mux2_1
X_10693_ VPWR VGND VPWR VGND _10692_/X _08195_/C _10693_/B1 _10693_/X sky130_fd_sc_hd__a21o_1
X_15220_ hold205/A _15220_/CLK _15220_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12432_ VGND VPWR VGND VPWR _12432_/X _12662_/A1 _12428_/X _12431_/X _12662_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_16_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12363_ VGND VPWR VPWR VGND _12363_/X _14956_/Q _12370_/S _14915_/Q sky130_fd_sc_hd__mux2_1
X_15151_ _15151_/Q _15151_/CLK _15151_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13706__823 VPWR VGND VPWR VGND _15046_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_11314_ VPWR VGND VGND VPWR _11355_/S _11347_/B _11340_/A sky130_fd_sc_hd__nor2_4
X_12294_ VGND VPWR VPWR VGND _12294_/X _14881_/Q _12701_/S _15417_/Q sky130_fd_sc_hd__mux2_1
X_15082_ _15082_/Q clkload37/A _15082_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_844 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11245_ VPWR VGND VPWR VGND _11244_/X _11245_/A1 _11243_/X _11245_/Y sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14124__1241 VPWR VGND VPWR VGND _15543_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_11176_ VGND VPWR VPWR VGND _11176_/X _11175_/X _11176_/S _11174_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13909__1026 VPWR VGND VPWR VGND _15281_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_10127_ VPWR VGND VPWR VGND _10126_/X _10616_/A1 _10125_/X _10127_/Y sky130_fd_sc_hd__a21oi_1
X_10058_ VPWR VGND VPWR VGND _12807_/B1 _10058_/A1 _12807_/A1 _15638_/D _10057_/Y
+ sky130_fd_sc_hd__a22o_1
X_14935_ hold922/A _14935_/CLK _14935_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14866_ hold993/A _14866_/CLK _14866_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14797_ hold732/A _14797_/CLK _14797_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15418_ hold786/A _15418_/CLK _15418_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15349_ _15349_/Q _15349_/CLK _15349_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13449__566 VPWR VGND VPWR VGND _14724_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
Xhold148 hold148/X hold148/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ VGND VPWR VPWR VGND _14140_/Q _09912_/A _09931_/B _09910_/X sky130_fd_sc_hd__or3b_1
Xhold159 hold159/X hold159/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout606 VPWR VGND _08405_/S _08408_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout639 VPWR VGND _09622_/S _09591_/Y VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout617 VGND VPWR _11441_/Y _11538_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09841_ VGND VPWR VPWR VGND _14181_/D hold470/X _09861_/S fanout69/X sky130_fd_sc_hd__mux2_1
Xfanout628 VPWR VGND _09756_/S _09729_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_09772_ VGND VPWR VPWR VGND _14277_/D fanout70/X _09792_/S hold575/X sky130_fd_sc_hd__mux2_1
XFILLER_39_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08723_ VGND VPWR VGND VPWR _15272_/D hold1009/X _08731_/A2 _08722_/X _11294_/A sky130_fd_sc_hd__o211a_1
XFILLER_73_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_54_512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_2_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08654_ VGND VPWR VGND VPWR _08714_/A2 _14381_/Q _08194_/B _08654_/X sky130_fd_sc_hd__o21ba_1
X_08585_ VPWR VGND VGND VPWR _15552_/Q _08585_/Y _09024_/A sky130_fd_sc_hd__nand2_1
X_07605_ VPWR VGND VPWR VGND _07908_/B1 _15636_/Q _07952_/A2 _07614_/A _11535_/A sky130_fd_sc_hd__a22o_1
X_07536_ VGND VPWR VPWR VGND _07536_/X _07535_/Y _07531_/A _07523_/Y _08591_/B _15561_/Q
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_14_Left_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07467_ VPWR VGND VGND VPWR _07468_/B _15449_/Q _07467_/B sky130_fd_sc_hd__or2_1
X_09206_ VGND VPWR VPWR VGND _14887_/D hold1068/X _09213_/S fanout67/X sky130_fd_sc_hd__mux2_1
X_07398_ VPWR VGND _07398_/X _07693_/B _07679_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_33_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09137_ VGND VPWR VPWR VGND _14961_/D fanout68/X _09157_/S hold738/X sky130_fd_sc_hd__mux2_1
X_09068_ VGND VPWR VPWR VGND _15025_/D hold1114/X _09090_/S fanout68/X sky130_fd_sc_hd__mux2_1
X_08019_ VPWR VGND VPWR VGND _07795_/C _07998_/B _07790_/B _08019_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_1384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold671 hold671/X hold671/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 hold660/X hold660/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ VGND VPWR VPWR VGND _11030_/X hold925/A _11175_/S hold469/A sky130_fd_sc_hd__mux2_1
Xhold693 hold693/X hold693/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 hold682/X hold682/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13242__359 VPWR VGND VPWR VGND _14517_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_79_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1360 hold1360/X _14925_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1393 hold1393/X _14129_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 hold1371/X _14137_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14720_ _14720_/Q _14720_/CLK _14720_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold1382 _09488_/A _14570_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11932_ VPWR VGND VGND VPWR _11932_/X hold678/A _12043_/B sky130_fd_sc_hd__or2_1
XFILLER_79_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14651_ hold679/A _14651_/CLK _14651_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11863_ VPWR VGND VGND VPWR _11844_/Y _11862_/X _10710_/B _15452_/Q _15452_/D _11296_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_707 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_60_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10814_ VPWR VGND VGND VPWR _10814_/X _10851_/A _10814_/B sky130_fd_sc_hd__or2_1
X_13095__212 VPWR VGND VPWR VGND _14338_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_11794_ VPWR VGND VGND VPWR _11794_/X _12591_/S _11794_/B sky130_fd_sc_hd__or2_1
X_14582_ hold668/A _14582_/CLK _14582_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10745_ VGND VPWR VGND VPWR _10745_/X _10742_/X _10744_/X _10745_/A1 _10745_/C1 sky130_fd_sc_hd__a211o_1
X_10676_ VGND VPWR VPWR VGND _10676_/X _14491_/Q _10696_/S hold683/A sky130_fd_sc_hd__mux2_1
X_13136__253 VPWR VGND VPWR VGND _14411_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_15203_ hold252/A _15203_/CLK _15203_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12415_ VGND VPWR VGND VPWR _12415_/X _12412_/X _12414_/X _12720_/A1 _12415_/C1 sky130_fd_sc_hd__a211o_1
X_12346_ VPWR VGND VGND VPWR _12346_/X hold405/A _12372_/S sky130_fd_sc_hd__or2_1
X_15134_ _15134_/Q _15134_/CLK _15134_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12277_ VGND VPWR VPWR VGND _12277_/X _12274_/X _12698_/S _12273_/X sky130_fd_sc_hd__mux2_1
X_15065_ _15065_/Q clkload14/A _15065_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13793__910 VPWR VGND VPWR VGND _15165_/CLK clkload23/A sky130_fd_sc_hd__inv_2
X_11228_ VPWR VGND VPWR VGND _11227_/X _07691_/X _12602_/B1 _11228_/X sky130_fd_sc_hd__a21o_1
X_11159_ VGND VPWR VPWR VGND _11159_/X hold580/A _11167_/S hold403/A sky130_fd_sc_hd__mux2_1
XFILLER_36_501 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13834__951 VPWR VGND VPWR VGND _15206_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
XFILLER_76_681 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_3_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14918_ hold382/A _14918_/CLK _14918_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14849_ _14849_/Q clkload20/A _14849_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08370_ VGND VPWR VPWR VGND _15403_/D hold734/X _08375_/S _09550_/A1 sky130_fd_sc_hd__mux2_1
X_07321_ VPWR VGND _07634_/B _07663_/B _07663_/A _07170_/Y _07320_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_07252_ VPWR VGND VGND VPWR _15457_/Q _07252_/B _08067_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_957 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_34_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_1362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07183_ VGND VPWR _07304_/A2 _07304_/B1 _07345_/C _14395_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_69_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout414 VGND VPWR fanout424/X _08178_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout403 VGND VPWR _10846_/A1 _11215_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout447 VPWR VGND _11210_/A _07691_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout436 VGND VPWR _11245_/A1 _11181_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout425 VGND VPWR _10634_/C1 _10608_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09824_ VGND VPWR VPWR VGND _14228_/D fanout7/X _09825_/S hold338/X sky130_fd_sc_hd__mux2_1
Xfanout469 VGND VPWR _12080_/A2 _12861_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout458 VPWR VGND _11246_/S _11209_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09755_ VGND VPWR VPWR VGND _14291_/D _09825_/A1 _09763_/S hold169/X sky130_fd_sc_hd__mux2_1
X_08706_ VGND VPWR VGND VPWR _08706_/X _08714_/A2 _08722_/C1 hold1453/X _08705_/X
+ sky130_fd_sc_hd__a211o_1
X_09686_ VGND VPWR VPWR VGND _14354_/D hold965/X _09693_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_13577__694 VPWR VGND VPWR VGND _14908_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_76_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08637_ VPWR VGND VPWR VGND hold1448/X _08700_/A2 _08637_/X _08662_/B1 _08636_/X
+ _08700_/B1 sky130_fd_sc_hd__a221o_1
XFILLER_74_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08568_ VPWR VGND VGND VPWR _08605_/A _08983_/B _08568_/Y sky130_fd_sc_hd__nor2_1
Xfanout10 VGND VPWR fanout9/A fanout10/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout21 VGND VPWR _08051_/X fanout21/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_08499_ VGND VPWR VPWR VGND _14138_/Q _14137_/Q _14139_/Q _09923_/D sky130_fd_sc_hd__or3_2
X_07519_ VGND VPWR _07519_/B _07519_/Y _15468_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
Xfanout43 VPWR VGND VGND VPWR clone6/A clone44/A sky130_fd_sc_hd__buf_8
Xfanout32 VGND VPWR fanout34/X fanout32/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout65 VGND VPWR fanout67/X fanout65/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout54 VPWR VGND VGND VPWR clone5/A fanout54/X sky130_fd_sc_hd__buf_8
XFILLER_50_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout87 VPWR VGND fanout87/X fanout88/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout98 VPWR VGND fanout98/X _08284_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_10530_ VPWR VGND VGND VPWR _10530_/X hold187/A _10627_/S sky130_fd_sc_hd__or2_1
X_13908__1025 VPWR VGND VPWR VGND _15280_/CLK clkload13/A sky130_fd_sc_hd__inv_2
Xfanout76 VPWR VGND VGND VPWR fanout79/X fanout76/X sky130_fd_sc_hd__buf_8
X_14123__1240 VPWR VGND VPWR VGND _15542_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_15265__940 _15265_/D _15265__940/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_10461_ VGND VPWR VPWR VGND _10465_/B hold879/A _10464_/S hold189/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12200_ VGND VPWR VPWR VGND _12200_/X hold584/A _12228_/B hold237/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10392_ VGND VPWR VGND VPWR _10392_/X _10698_/A1 _10388_/X _10391_/X _10697_/B1 sky130_fd_sc_hd__o211a_1
X_12131_ VGND VPWR VPWR VGND _12135_/B hold721/A _12155_/S hold159/A sky130_fd_sc_hd__mux2_1
XFILLER_2_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold490 hold490/X hold490/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12062_ VGND VPWR VGND VPWR _12062_/X _12230_/A1 _12058_/X _12061_/X _12226_/C1 sky130_fd_sc_hd__o211a_1
X_11013_ VGND VPWR VGND VPWR _11013_/X _11185_/A1 _11009_/X _11012_/X _11185_/C1 sky130_fd_sc_hd__o211a_1
X_13818__935 VPWR VGND VPWR VGND _15190_/CLK clkload48/A sky130_fd_sc_hd__inv_2
Xhold1190 hold1190/X _15339_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14703_ hold675/A _14703_/CLK _14703_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_545 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11915_ VGND VPWR VPWR VGND _11915_/X _11912_/X _12069_/S _11911_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_824 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_526 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_57_1362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11846_ VGND VPWR VPWR VGND _11846_/X hold965/A _12089_/S hold583/A sky130_fd_sc_hd__mux2_1
X_14634_ _14634_/Q _14634_/CLK _14634_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14565_ hold695/A _14565_/CLK _14565_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11777_ VGND VPWR VGND VPWR _11777_/X _11776_/X _11775_/X _12106_/S _12017_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_18_1357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13370__487 VPWR VGND VPWR VGND _14645_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_10728_ VGND VPWR VPWR VGND _10729_/B _10727_/Y _10728_/S _10719_/Y sky130_fd_sc_hd__mux2_1
X_14496_ _14496_/Q _14496_/CLK _14496_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkload24 VGND VPWR VGND VPWR clkload24/A clkload24/Y sky130_fd_sc_hd__clkinv_8
Xclkload13 VGND VPWR VPWR VGND clkload13/A clkload13/Y sky130_fd_sc_hd__clkinv_2
X_10659_ VGND VPWR VGND VPWR _10659_/X _10658_/X _10657_/X _10557_/A _10717_/C1 sky130_fd_sc_hd__a211o_1
Xclkload35 clkload35/Y clkload35/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload46 VGND VPWR VGND VPWR clkload46/Y clkload46/A sky130_fd_sc_hd__inv_12
X_12329_ VPWR VGND VGND VPWR _12329_/X hold387/A _12339_/B sky130_fd_sc_hd__or2_1
X_15117_ hold985/A _15117_/CLK _15117_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15048_ hold595/A _15048_/CLK _15048_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07870_ VGND VPWR VPWR VGND _07870_/D _07870_/C _07870_/B _07870_/A clone5/A sky130_fd_sc_hd__or4_4
X_13264__381 VPWR VGND VPWR VGND _14539_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
XFILLER_37_810 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09540_ VGND VPWR VPWR VGND _14522_/D fanout28/X _09555_/S hold241/X sky130_fd_sc_hd__mux2_1
XFILLER_37_876 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09471_ VGND VPWR VPWR VGND _14585_/D fanout24/X _09485_/S hold245/X sky130_fd_sc_hd__mux2_1
X_08422_ VPWR VGND VGND VPWR _14128_/Q _14126_/Q _08422_/C _08425_/A sky130_fd_sc_hd__nor3_2
X_13611__728 VPWR VGND VPWR VGND _14951_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_08353_ VGND VPWR VPWR VGND _15420_/D hold590/X _08372_/S clone5/X sky130_fd_sc_hd__mux2_1
X_07304_ VPWR VGND VGND VPWR _14399_/Q _07304_/A2 _07304_/B1 _07306_/B sky130_fd_sc_hd__o21a_1
X_08284_ VGND VPWR VGND VPWR _08299_/A2 _15607_/Q _08283_/X _08284_/X sky130_fd_sc_hd__a21o_2
XFILLER_50_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07235_ VPWR VGND VPWR VGND _10062_/A _08239_/A _07219_/X _08222_/B sky130_fd_sc_hd__a21o_1
Xclkload7 VGND VPWR VPWR VGND clkload7/A clkload7/Y sky130_fd_sc_hd__clkinv_2
X_07166_ VPWR VGND VGND VPWR _15472_/Q _07166_/B _07338_/B sky130_fd_sc_hd__nor2_1
X_07097_ VPWR VGND VPWR VGND _07222_/B _15447_/Q sky130_fd_sc_hd__inv_2
X_13505__622 VPWR VGND VPWR VGND _14780_/CLK clkload20/A sky130_fd_sc_hd__inv_2
Xfanout222 VGND VPWR fanout234/X _12189_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout200 VGND VPWR _11894_/S _11958_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout211 VGND VPWR _12674_/A1 _12670_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout233 VPWR VGND _12572_/C1 fanout234/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout255 VPWR VGND _12864_/A1 _07936_/X VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_43_1417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout244 VPWR VGND _12415_/C1 _12376_/B2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout277 VPWR VGND _12866_/A1 fanout282/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout266 VPWR VGND _12214_/A _07912_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout299 VGND VPWR _10484_/B _10169_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07999_ VPWR VGND VGND VPWR _07999_/X _07999_/A _07999_/B sky130_fd_sc_hd__or2_1
Xfanout288 VGND VPWR _10140_/S _10604_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09807_ VGND VPWR VPWR VGND _14245_/D fanout70/X _09827_/S hold283/X sky130_fd_sc_hd__mux2_1
X_09738_ VGND VPWR VPWR VGND _14308_/D fanout66/X _09757_/S hold370/X sky130_fd_sc_hd__mux2_1
X_09669_ VGND VPWR VPWR VGND _14371_/D hold776/X _09690_/S fanout62/X sky130_fd_sc_hd__mux2_1
X_12680_ VGND VPWR VPWR VGND _12680_/X hold513/A _12689_/S hold553/A sky130_fd_sc_hd__mux2_1
X_11700_ VPWR VGND VGND VPWR _11700_/X hold499/A _12052_/S sky130_fd_sc_hd__or2_1
XFILLER_39_1070 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11631_ VPWR VGND VGND VPWR _11631_/X hold233/A _12117_/B sky130_fd_sc_hd__or2_1
X_11562_ VPWR VGND VPWR VGND _11561_/Y _11563_/B _11542_/A _15441_/D sky130_fd_sc_hd__a21oi_1
X_14350_ _14350_/Q _14350_/CLK _14350_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_24_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10513_ VGND VPWR VPWR VGND _10513_/X hold994/A _10520_/S hold650/A sky130_fd_sc_hd__mux2_1
XFILLER_10_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14281_ hold557/A _14281_/CLK _14281_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11493_ VGND VPWR VPWR VGND _11493_/X _15083_/Q _11535_/C _15081_/Q sky130_fd_sc_hd__mux2_1
X_10444_ VPWR VGND VGND VPWR _10444_/X _10662_/S _10444_/B sky130_fd_sc_hd__or2_1
X_10375_ VGND VPWR VGND VPWR _10375_/X _10372_/X _10374_/X _10698_/A1 _10693_/B1 sky130_fd_sc_hd__a211o_1
X_13248__365 VPWR VGND VPWR VGND _14523_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_12114_ VGND VPWR VGND VPWR _12114_/X hold917/A _12118_/A2 _12118_/B1 _12113_/X sky130_fd_sc_hd__o211a_1
XFILLER_3_975 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12045_ VGND VPWR VGND VPWR _12045_/X _12042_/X _12044_/X _12156_/A1 _12212_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_59_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12878_ VPWR VGND VPWR VGND _12878_/B _12878_/C _12878_/A _12878_/X _08197_/S sky130_fd_sc_hd__or4b_1
X_11829_ VGND VPWR VPWR VGND _11829_/X hold761/A _12183_/S hold265/A sky130_fd_sc_hd__mux2_1
X_14617_ hold521/A _14617_/CLK _14617_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15597_ _15597_/Q clkload55/A _15597_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14548_ hold455/A _14548_/CLK _14548_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14479_ hold968/A _14479_/CLK _14479_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08971_ VGND VPWR VPWR VGND _08972_/B _07560_/D _09906_/A hold758/A sky130_fd_sc_hd__mux2_1
X_07922_ VGND VPWR _07922_/B _07923_/B _07925_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_69_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_64_1196 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07853_ VGND VPWR VGND VPWR _10891_/C1 _08286_/A _07870_/C _07914_/B1 sky130_fd_sc_hd__a21oi_2
X_13907__1024 VPWR VGND VPWR VGND _15279_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_07784_ VPWR VGND VPWR VGND _07783_/B _08126_/A _07747_/X _08097_/A sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09523_ VPWR VGND VGND VPWR _09523_/X _09523_/A _09549_/S sky130_fd_sc_hd__or2_1
X_13041__158 VPWR VGND VPWR VGND _14284_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_52_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09454_ _14602_/D fanout94/X fanout90/X _09452_/Y _09453_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08405_ VGND VPWR VPWR VGND _15372_/D _09792_/A1 _08405_/S hold398/X sky130_fd_sc_hd__mux2_1
X_09385_ VGND VPWR VPWR VGND _09408_/S hold1096/X fanout81/X _14664_/D sky130_fd_sc_hd__mux2_2
XFILLER_75_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08336_ VGND VPWR VPWR VGND _15483_/D _09691_/A0 _08338_/S hold809/X sky130_fd_sc_hd__mux2_1
X_08267_ VGND VPWR VPWR VGND _15515_/D _09691_/A0 _08267_/S hold355/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_67_Right_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08198_ VGND VPWR VPWR VGND _08198_/X _08197_/X _08198_/S _08196_/X sky130_fd_sc_hd__mux2_1
X_07218_ VGND VPWR VPWR VGND _07234_/B _07220_/S _15593_/Q _14382_/Q sky130_fd_sc_hd__mux2_4
X_07149_ VPWR VGND _07411_/A _07149_/B _15476_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_10160_ VPWR VGND VGND VPWR _10160_/X hold215/A _10464_/S sky130_fd_sc_hd__or2_1
X_10091_ VGND VPWR VPWR VGND _10095_/B hold611/A _10602_/S hold320/A sky130_fd_sc_hd__mux2_1
XFILLER_43_1247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Right_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12801_ VPWR VGND VGND VPWR _12822_/A _08005_/Y _10056_/A _12801_/X sky130_fd_sc_hd__o21a_1
X_10993_ VGND VPWR VPWR VGND _10993_/X hold939/A _10994_/S hold754/A sky130_fd_sc_hd__mux2_1
X_13633__750 VPWR VGND VPWR VGND _14973_/CLK clkload49/A sky130_fd_sc_hd__inv_2
X_15520_ hold447/A _15520_/CLK _15520_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12732_ VPWR VGND VGND VPWR _12732_/A _12732_/B _12732_/Y sky130_fd_sc_hd__nor2_1
X_15451_ _15451_/Q clkload55/A _15451_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_15_378 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14402_ _14402_/Q clkload41/A _14402_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12663_ VGND VPWR VPWR VGND _12663_/X _14440_/Q _12664_/S _14696_/Q sky130_fd_sc_hd__mux2_1
X_12594_ VPWR VGND VGND VPWR _12594_/X _14994_/Q _12594_/B sky130_fd_sc_hd__or2_1
X_15382_ hold528/A _15382_/CLK _15382_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11614_ VGND VPWR VPWR VGND _11614_/X hold512/A _11838_/S hold541/A sky130_fd_sc_hd__mux2_1
XFILLER_7_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_1305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11545_ VPWR VGND VGND VPWR _11545_/A _11545_/Y _11545_/B sky130_fd_sc_hd__nand2_1
X_14333_ hold690/A _14333_/CLK _14333_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_522 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11476_ VGND VPWR VPWR VGND _11476_/X _11475_/X _11476_/S _15456_/Q sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Left_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14264_ hold383/A _14264_/CLK _14264_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10427_ VGND VPWR VPWR VGND _10427_/X hold357/A _10742_/S hold338/A sky130_fd_sc_hd__mux2_1
X_14195_ _14195_/Q _14195_/CLK _14195_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13482__599 VPWR VGND VPWR VGND _14757_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_10358_ VGND VPWR VPWR VGND _10359_/B _10357_/Y _10617_/S _10349_/Y sky130_fd_sc_hd__mux2_1
X_10289_ VPWR VGND VGND VPWR _10289_/X hold362/A _10521_/B sky130_fd_sc_hd__or2_1
XFILLER_78_551 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12028_ VGND VPWR VPWR VGND _12029_/B _12027_/Y _12102_/S _12019_/Y sky130_fd_sc_hd__mux2_1
X_14102__1219 VPWR VGND VPWR VGND _15521_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_59_1210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_695 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13376__493 VPWR VGND VPWR VGND _14651_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_72_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09170_ VGND VPWR VPWR VGND _14921_/D hold354/X _09194_/S fanout73/X sky130_fd_sc_hd__mux2_1
X_08121_ VPWR VGND VPWR VGND _08293_/A3 _15074_/Q _11440_/B _08121_/X _07241_/X sky130_fd_sc_hd__a22o_1
X_08052_ VGND VPWR VPWR VGND _15526_/D fanout21/X _08267_/S hold238/X sky130_fd_sc_hd__mux2_1
XFILLER_0_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08954_ VPWR VGND VPWR VGND _08969_/A hold1428/X _08933_/A _08954_/X _15119_/Q sky130_fd_sc_hd__a22o_1
X_07905_ VPWR VGND VGND VPWR _15563_/Q _07931_/A _07906_/B sky130_fd_sc_hd__nor2_1
X_08885_ VGND VPWR VGND VPWR _15150_/D hold1294/X _08919_/A2 _08884_/X _11388_/S sky130_fd_sc_hd__o211a_1
X_07836_ VGND VPWR _08022_/B _15555_/Q _15556_/Q _08059_/B VPWR VGND sky130_fd_sc_hd__and3_1
X_07767_ VPWR VGND VPWR VGND _07826_/D _15591_/Q _07765_/B _08272_/B _09164_/A sky130_fd_sc_hd__a22o_1
X_13617__734 VPWR VGND VPWR VGND _14957_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_09506_ VGND VPWR VPWR VGND _14553_/D fanout24/X _09520_/S hold1018/X sky130_fd_sc_hd__mux2_1
X_07698_ VGND VPWR VGND VPWR _07698_/X _07881_/A2 _07696_/X _15089_/Q _07697_/X sky130_fd_sc_hd__a211o_1
X_09437_ VGND VPWR VPWR VGND _14615_/D fanout15/X _09449_/S hold547/X sky130_fd_sc_hd__mux2_1
X_14199__917 _14199_/D _14199__917/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09368_ VGND VPWR VPWR VGND _14678_/D hold815/X _09379_/S fanout12/X sky130_fd_sc_hd__mux2_1
XFILLER_24_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08319_ VGND VPWR VPWR VGND _15500_/D fanout41/X _08332_/S hold881/X sky130_fd_sc_hd__mux2_1
X_09299_ VGND VPWR VPWR VGND _14742_/D fanout12/X _09310_/S hold284/X sky130_fd_sc_hd__mux2_1
X_11330_ VPWR VGND _11330_/X _11408_/A _14829_/Q _14833_/Q _11340_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XANTENNA_82 _08190_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_71 _09864_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_60 fanout539/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_93 _14406_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11261_ VPWR VGND VGND VPWR _11261_/X _14998_/Q _11261_/B sky130_fd_sc_hd__or2_1
X_10212_ VGND VPWR VPWR VGND _10212_/X hold833/A _10567_/S hold672/A sky130_fd_sc_hd__mux2_1
X_11192_ VPWR VGND VGND VPWR _11173_/Y _11191_/X _12677_/A2 _14408_/Q _14408_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_10143_ VGND VPWR VPWR VGND _10143_/X hold871/A _10604_/S hold648/A sky130_fd_sc_hd__mux2_1
XFILLER_75_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10074_ VGND VPWR VPWR VGND _10074_/X _10074_/A1 _10074_/S _10074_/A0 sky130_fd_sc_hd__mux2_1
X_14951_ hold992/A _14951_/CLK _14951_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14882_ hold846/A _14882_/CLK _14882_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_36_908 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13063__180 VPWR VGND VPWR VGND _14306_/CLK clkload42/A sky130_fd_sc_hd__inv_2
XFILLER_78_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10976_ VGND VPWR VGND VPWR _10976_/X _11004_/A1 _10972_/X _10975_/X _11235_/C1 sky130_fd_sc_hd__o211a_1
X_15503_ _15503_/Q _15503_/CLK _15503_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_43_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12715_ VGND VPWR VPWR VGND _12719_/B _14634_/Q _12726_/S _14666_/Q sky130_fd_sc_hd__mux2_1
X_15434_ _15434_/Q clkload47/A _15434_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12646_ VGND VPWR VGND VPWR _12646_/X _12662_/A1 _12642_/X _12645_/X _12662_/C1 sky130_fd_sc_hd__o211a_1
X_15365_ _15365_/Q _15365_/CLK hold154/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13410__527 VPWR VGND VPWR VGND _14685_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_12577_ VGND VPWR VPWR VGND _12577_/X _14214_/Q _12577_/S _15222_/Q sky130_fd_sc_hd__mux2_1
X_13906__1023 VPWR VGND VPWR VGND _15278_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_14316_ hold780/A _14316_/CLK _14316_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold308 hold308/X hold308/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11528_ VGND VPWR VPWR VGND _15093_/D _11527_/X _11528_/S hold1394/X sky130_fd_sc_hd__mux2_1
X_15296_ hold907/A _15296_/CLK _15296_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11459_ VGND VPWR VPWR VGND _15070_/D _11458_/X _11480_/S hold1386/X sky130_fd_sc_hd__mux2_1
X_14247_ _14247_/Q _14247_/CLK _14247_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold319 hold319/X hold319/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14178_ hold825/A _14178_/CLK _14178_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13304__421 VPWR VGND VPWR VGND _14579_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
Xhold1008 hold1008/X _15284_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 hold1019/X _14476_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08670_ VPWR VGND VPWR VGND _15290_/Q _08562_/A _08670_/X _08691_/B1 _08669_/X _08700_/B1
+ sky130_fd_sc_hd__a221o_1
X_07621_ VPWR VGND VGND VPWR _07637_/A _07621_/B _07625_/A _07621_/Y sky130_fd_sc_hd__nor3_1
X_07552_ VGND VPWR VPWR VGND _07560_/D _07551_/X _07523_/Y _07500_/Y _07552_/B1 _15559_/Q
+ sky130_fd_sc_hd__a32o_1
X_14082__1199 VPWR VGND VPWR VGND _15501_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_07483_ VPWR VGND VGND VPWR _07483_/A _07580_/B _07483_/B sky130_fd_sc_hd__nand2_1
X_09222_ VGND VPWR VPWR VGND _14871_/D hold1051/X _09229_/S fanout5/X sky130_fd_sc_hd__mux2_1
X_09153_ VGND VPWR VPWR VGND _14945_/D fanout8/X _09163_/S hold830/X sky130_fd_sc_hd__mux2_1
XFILLER_33_1224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_679 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08104_ VPWR VGND VGND VPWR _08104_/A _08104_/B _08104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09084_ VGND VPWR VPWR VGND _15009_/D hold1004/X _09094_/S fanout10/X sky130_fd_sc_hd__mux2_1
X_08035_ VGND VPWR VPWR VGND _08035_/X _08034_/X _08195_/A _07616_/X sky130_fd_sc_hd__mux2_1
Xhold820 hold820/X hold820/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 hold853/X hold853/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 hold842/X hold842/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 hold831/X hold831/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 hold864/X hold864/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 hold886/X hold886/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_1017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold897 hold897/X hold897/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 hold875/X hold875/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ VPWR VGND VGND VPWR _15609_/Q _09986_/B _09987_/B sky130_fd_sc_hd__nor2_1
X_08937_ VGND VPWR _09869_/A _09873_/A _08937_/Y _15479_/Q VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_44_1364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13047__164 VPWR VGND VPWR VGND _14290_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_08868_ VPWR VGND VGND VPWR _08868_/X _15158_/Q _08868_/B sky130_fd_sc_hd__or2_1
XFILLER_79_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07819_ VPWR VGND VGND VPWR _07819_/A _07820_/B _07856_/A sky130_fd_sc_hd__nand2_1
X_08799_ VGND VPWR VPWR VGND _15210_/D fanout27/X _08806_/S hold328/X sky130_fd_sc_hd__mux2_1
X_13851__968 VPWR VGND VPWR VGND _15223_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_10830_ VGND VPWR VGND VPWR _10830_/X _11096_/C1 _10825_/X _10829_/X _11218_/C1 sky130_fd_sc_hd__o211a_1
X_10761_ VPWR VGND VGND VPWR _10761_/X _11092_/S _10761_/B sky130_fd_sc_hd__or2_1
XFILLER_13_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10692_ VGND VPWR VPWR VGND _10692_/X _14363_/Q _10702_/S hold409/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12500_ VPWR VGND VPWR VGND _12499_/X _12656_/A1 _12498_/X _12500_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12431_ VPWR VGND VGND VPWR _12431_/X _12655_/S _12431_/B sky130_fd_sc_hd__or2_1
X_13745__862 VPWR VGND VPWR VGND _15117_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_12362_ VGND VPWR VPWR VGND _12365_/B _14368_/Q _12599_/S _14720_/Q sky130_fd_sc_hd__mux2_1
X_15150_ _15150_/Q _15150_/CLK _15150_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14101__1218 VPWR VGND VPWR VGND _15520_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_11313_ VPWR VGND VGND VPWR _14822_/Q _11421_/A _11347_/B _11313_/C sky130_fd_sc_hd__nand3_1
X_12293_ VGND VPWR VGND VPWR _12293_/X hold743/A _12705_/A2 _12256_/S _12292_/X sky130_fd_sc_hd__o211a_1
X_15081_ _15081_/Q clkload37/A _15081_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11244_ VGND VPWR VPWR VGND _11244_/X _11241_/X _11244_/S _11240_/X sky130_fd_sc_hd__mux2_1
X_11175_ VGND VPWR VPWR VGND _11175_/X _14376_/Q _11175_/S _14728_/Q sky130_fd_sc_hd__mux2_1
XFILLER_62_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10126_ VGND VPWR VPWR VGND _10126_/X _10123_/X _10615_/S _10122_/X sky130_fd_sc_hd__mux2_1
X_14934_ _14934_/Q clkload29/A _14934_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10057_ VPWR VGND VGND VPWR _14803_/Q _14801_/Q _10057_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14865_ _14865_/Q _14865_/CLK _14865_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_63_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14796_ _14796_/Q _14796_/CLK _14796_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10959_ VGND VPWR VGND VPWR _10959_/X _11181_/A1 _10954_/X _10958_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_32_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15417_ _15417_/Q _15417_/CLK _15417_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12629_ VGND VPWR VGND VPWR _12629_/X _12740_/A1 _12624_/X _12628_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_15348_ _15348_/Q _15348_/CLK _15348_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15279_ _15279_/Q _15279_/CLK _15279_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold149 hold149/X hold149/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_1326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09840_ VGND VPWR VPWR VGND _14182_/D _09861_/S hold1123/X fanout74/X sky130_fd_sc_hd__mux2_4
Xfanout629 _09757_/S _09760_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout607 VPWR VGND _08393_/S _08408_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout618 VGND VPWR _11441_/Y _11528_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09771_ VGND VPWR VPWR VGND _14278_/D _09795_/S clone47/A hold1260/X sky130_fd_sc_hd__mux2_4
XFILLER_67_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08722_ VPWR VGND VPWR VGND hold976/A _08523_/B _08722_/X _08728_/B1 _14383_/Q _08722_/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08653_ VGND VPWR VGND VPWR _15295_/D hold1046/X _08721_/A2 _08652_/X _11937_/C1
+ sky130_fd_sc_hd__o211a_1
X_08584_ VGND VPWR VGND VPWR _15310_/D hold990/X _08613_/A2 _08583_/X _09000_/C1 sky130_fd_sc_hd__o211a_1
X_07604_ VGND VPWR VGND VPWR _07914_/B1 _07418_/B _07603_/X _07614_/B sky130_fd_sc_hd__o21ba_1
X_07535_ VGND VPWR _07530_/A _07530_/C _07535_/Y _07530_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
X_13688__805 VPWR VGND VPWR VGND _15028_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_07466_ VPWR VGND VGND VPWR _15449_/Q _07487_/A _07467_/B sky130_fd_sc_hd__nand2_1
X_09205_ VGND VPWR VPWR VGND _14888_/D hold935/X _09213_/S fanout69/X sky130_fd_sc_hd__mux2_1
X_13729__846 VPWR VGND VPWR VGND _15101_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_07397_ VPWR VGND VPWR VGND _07397_/B _07397_/C _07397_/A _07694_/B sky130_fd_sc_hd__or3_1
XFILLER_33_1021 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09136_ VGND VPWR VPWR VGND _14962_/D fanout73/X _09160_/S hold458/X sky130_fd_sc_hd__mux2_1
X_09067_ VGND VPWR VPWR VGND _15026_/D _09088_/S hold1268/X clone111/X sky130_fd_sc_hd__mux2_4
X_08018_ VPWR VGND VGND VPWR _08017_/X _07421_/Y _08016_/X _07421_/A _08032_/B _07996_/X
+ sky130_fd_sc_hd__o221a_1
Xhold661 hold661/X hold661/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 hold650/X hold650/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1396 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold672 hold672/X hold672/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold683 hold683/X hold683/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 hold694/X hold694/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ VGND VPWR VGND VPWR _09969_/X _09970_/A _08862_/C _15480_/Q _09024_/A sky130_fd_sc_hd__o211a_1
X_13281__398 VPWR VGND VPWR VGND _14556_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
XFILLER_79_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1350 _09988_/A _15610_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1361 hold1361/X _15069_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1383 hold1383/X _14127_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13905__1022 VPWR VGND VPWR VGND _15277_/CLK clkload14/A sky130_fd_sc_hd__inv_2
Xhold1372 hold1372/X _14698_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 hold1394/X _15093_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11931_ VGND VPWR VPWR VGND _11931_/X hold812/A _12043_/B hold696/A sky130_fd_sc_hd__mux2_1
X_11862_ VPWR VGND VPWR VGND _11861_/X _12103_/A _12121_/B1 _11862_/X sky130_fd_sc_hd__a21o_1
X_14650_ hold676/A _14650_/CLK _14650_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14581_ hold497/A _14581_/CLK _14581_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10813_ VGND VPWR VPWR VGND _10813_/X hold568/A _11223_/S hold261/A sky130_fd_sc_hd__mux2_1
X_11793_ VGND VPWR VPWR VGND _11793_/X _14545_/Q _12589_/S hold349/A sky130_fd_sc_hd__mux2_1
X_13175__292 VPWR VGND VPWR VGND _14450_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_10744_ VGND VPWR VGND VPWR _10744_/X _15016_/Q _10744_/A2 _10743_/X _10732_/S sky130_fd_sc_hd__o211a_1
X_10675_ VGND VPWR VPWR VGND _10675_/X hold639/A _10696_/S hold679/A sky130_fd_sc_hd__mux2_1
XFILLER_9_458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15202_ hold225/A _15202_/CLK _15202_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12414_ VGND VPWR VGND VPWR _12414_/X _15021_/Q _12488_/A2 _12721_/S _12413_/X sky130_fd_sc_hd__o211a_1
X_12345_ VGND VPWR VPWR VGND _12345_/X _14624_/Q _12372_/S hold379/A sky130_fd_sc_hd__mux2_1
XFILLER_64_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15133_ _15133_/Q _15133_/CLK _15133_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12974__91 VPWR VGND VPWR VGND _14217_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_15064_ _15697_/A _15064_/CLK _15064_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12276_ VGND VPWR VGND VPWR _12276_/X _12256_/S _12272_/X _12275_/X _12702_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_4_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14081__1198 VPWR VGND VPWR VGND _15500_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_11227_ VPWR VGND _11227_/X _11226_/X _11222_/X _10765_/S _11218_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_13522__639 VPWR VGND VPWR VGND _14797_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_11158_ VGND VPWR VPWR VGND _11158_/X _14344_/Q _11167_/S hold247/A sky130_fd_sc_hd__mux2_1
X_10109_ VGND VPWR VPWR VGND _10109_/X hold931/A _10516_/S hold192/A sky130_fd_sc_hd__mux2_1
X_11089_ VGND VPWR VGND VPWR _11089_/X _11096_/C1 _11084_/X _11088_/X _11218_/C1 sky130_fd_sc_hd__o211a_1
X_13873__990 VPWR VGND VPWR VGND _15245_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
XFILLER_48_384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14917_ hold834/A _14917_/CLK _14917_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1289 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14848_ _14848_/Q clkload20/A _14848_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1041 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07320_ VGND VPWR VGND VPWR _07338_/A _07338_/B _07339_/B _07320_/X sky130_fd_sc_hd__o21ba_1
X_14779_ hold601/A _14779_/CLK _14779_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13416__533 VPWR VGND VPWR VGND _14691_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XFILLER_34_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07251_ VPWR VGND _08041_/A _07252_/B _15457_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07182_ VPWR VGND VPWR VGND _07971_/A _07182_/A _07972_/A sky130_fd_sc_hd__or2_2
XFILLER_69_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout404 VGND VPWR _10846_/A1 _11086_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout448 VPWR VGND VGND VPWR _07690_/Y _10893_/B1 sky130_fd_sc_hd__buf_8
X_09823_ VGND VPWR VPWR VGND _14229_/D fanout8/X _09833_/S hold189/X sky130_fd_sc_hd__mux2_1
X_12983__100 VPWR VGND VPWR VGND _14226_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
Xfanout426 VGND VPWR _10634_/C1 _10616_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout437 VGND VPWR _11023_/A1 _11245_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout415 VGND VPWR _12868_/A1 _11235_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout459 VPWR VGND _10765_/S _11209_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09754_ VGND VPWR VPWR VGND _14292_/D fanout7/X _09756_/S hold292/X sky130_fd_sc_hd__mux2_1
X_14100__1217 VPWR VGND VPWR VGND _15519_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_09685_ VGND VPWR VPWR VGND _14355_/D hold861/X _09693_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
X_08705_ VGND VPWR VGND VPWR _08705_/X _14390_/Q _08664_/B _08711_/B1 _08649_/X sky130_fd_sc_hd__o211a_1
X_08636_ VPWR VGND VGND VPWR _08635_/X _08690_/S _08194_/Y _14409_/Q _08636_/X _08634_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_74_1143 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08567_ _08983_/B _08604_/B2 _08544_/B _08566_/X _08565_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xfanout11 VGND VPWR _08108_/X fanout9/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_13159__276 VPWR VGND VPWR VGND _14434_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_08498_ VPWR VGND VPWR VGND _08498_/Y _08500_/C sky130_fd_sc_hd__inv_2
X_07518_ VPWR VGND VPWR VGND _07539_/C _07539_/B _07539_/A _07518_/X sky130_fd_sc_hd__a21o_1
Xfanout44 VGND VPWR fanout45/X fanout44/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout33 VGND VPWR fanout34/X fanout33/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_74_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07449_ VPWR VGND VGND VPWR _15455_/Q _11535_/A _07450_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout66 VGND VPWR fanout67/X fanout66/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout88 VPWR VGND fanout88/X fanout89/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout99 VPWR VGND VPWR VGND fanout99/X _08284_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout77 VPWR VGND fanout77/X fanout79/X VPWR VGND sky130_fd_sc_hd__buf_6
X_10460_ VPWR VGND VPWR VGND _10459_/X _10706_/C1 _10458_/X _10460_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09119_ VGND VPWR VPWR VGND _14976_/D hold678/X _09126_/S fanout5/X sky130_fd_sc_hd__mux2_1
X_10391_ VPWR VGND VGND VPWR _10391_/X _10685_/S _10391_/B sky130_fd_sc_hd__or2_1
X_12130_ VPWR VGND VPWR VGND _12129_/X _12212_/A1 _12128_/X _12130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_1171 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12061_ VPWR VGND VGND VPWR _12061_/X _12221_/S _12061_/B sky130_fd_sc_hd__or2_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold480 hold480/X hold480/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold491 hold491/X hold491/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ VPWR VGND VGND VPWR _11012_/X _11176_/S _11012_/B sky130_fd_sc_hd__or2_1
X_13857__974 VPWR VGND VPWR VGND _15229_/CLK clkload24/A sky130_fd_sc_hd__inv_2
XFILLER_38_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13103__220 VPWR VGND VPWR VGND _14346_/CLK clkload33/A sky130_fd_sc_hd__inv_2
XFILLER_20_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1180 hold1180/X _14247_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14702_ hold468/A _14702_/CLK _14702_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold1191 hold1191/X _14632_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ VGND VPWR VGND VPWR _11914_/X _12230_/A1 _11910_/X _11913_/X _12202_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_46_899 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14633_ hold500/A _14633_/CLK _14633_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11845_ VGND VPWR VPWR VGND _11845_/X hold919/A _12117_/B hold435/A sky130_fd_sc_hd__mux2_1
XFILLER_57_1374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14564_ hold740/A _14564_/CLK _14564_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11776_ VGND VPWR VPWR VGND _11776_/X hold778/A _12006_/B hold734/A sky130_fd_sc_hd__mux2_1
X_14495_ hold847/A _14495_/CLK _14495_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10727_ VPWR VGND VPWR VGND _10726_/X _10745_/C1 _10725_/X _10727_/Y sky130_fd_sc_hd__a21oi_1
Xclkload25 VGND VPWR VGND VPWR clkload25/A clkload25/Y sky130_fd_sc_hd__bufinv_8
Xclkload14 clkload14/Y clkload14/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
X_10658_ VGND VPWR VPWR VGND _10658_/X hold828/A _10670_/S hold576/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1093 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkload47 VGND VPWR VGND VPWR clkload47/Y clkload47/A sky130_fd_sc_hd__inv_12
Xclkload36 VPWR VGND VPWR VGND clkload36/Y clkload36/A sky130_fd_sc_hd__inv_6
X_10589_ VGND VPWR VGND VPWR _10589_/X _10745_/C1 _10588_/X _10585_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_15116_ hold588/A _15116_/CLK _15116_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12328_ VGND VPWR VPWR VGND _12328_/X _12327_/X _12328_/S _12326_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12259_ VGND VPWR VPWR VGND _12259_/X hold979/A _12339_/B hold685/A sky130_fd_sc_hd__mux2_1
X_15047_ hold420/A _15047_/CLK _15047_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09470_ VGND VPWR VPWR VGND _14586_/D fanout29/X _09478_/S hold218/X sky130_fd_sc_hd__mux2_1
X_08421_ VPWR VGND VPWR VGND _14129_/Q _14127_/Q _14130_/Q _08422_/C sky130_fd_sc_hd__or3_1
XFILLER_51_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13650__767 VPWR VGND VPWR VGND _14990_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_12888__5 VPWR VGND VPWR VGND _14130_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08352_ VGND VPWR VPWR VGND _15421_/D hold425/X _08356_/S fanout56/X sky130_fd_sc_hd__mux2_1
X_08283_ VGND VPWR VGND VPWR _08283_/X _08271_/Y _08281_/X _10058_/A1 _08282_/X sky130_fd_sc_hd__a211o_1
X_07303_ VPWR VGND VGND VPWR _07876_/A _07813_/A _07311_/A sky130_fd_sc_hd__or2_1
X_07234_ VGND VPWR VGND VPWR _10062_/A _07234_/B _07234_/A sky130_fd_sc_hd__xnor2_4
Xclkload8 VGND VPWR VGND VPWR clkload8/Y clkload8/A sky130_fd_sc_hd__inv_12
X_07165_ VPWR VGND _07338_/A _07166_/B _15472_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_13904__1021 VPWR VGND VPWR VGND _15276_/CLK clkload14/A sky130_fd_sc_hd__inv_2
X_07096_ VPWR VGND VPWR VGND _07234_/A _15448_/Q sky130_fd_sc_hd__inv_2
X_13544__661 VPWR VGND VPWR VGND _14875_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
Xfanout201 VPWR VGND _11968_/S _11894_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout212 VGND VPWR fanout217/X _12674_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout223 VGND VPWR fanout234/X _12202_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout245 VPWR VGND _12376_/B2 _07955_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout234 fanout234/X _07956_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_43_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout256 VPWR VGND _12102_/S _12176_/S VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_75_906 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09806_ VGND VPWR VPWR VGND _14246_/D _09830_/S clone47/X hold1154/X sky130_fd_sc_hd__mux2_4
X_07998_ _07798_/A _07998_/B _07999_/B _07998_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
Xfanout278 VGND VPWR _11184_/A2 _11252_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout289 VGND VPWR fanout314/X _10140_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout267 VGND VPWR _12732_/A _12658_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09737_ VGND VPWR VPWR VGND _14309_/D fanout70/X _09757_/S hold373/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_66_clk clkload11/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09668_ VGND VPWR VPWR VGND _14372_/D hold955/X _09687_/S fanout67/X sky130_fd_sc_hd__mux2_1
X_08619_ VGND VPWR VGND VPWR _15303_/D hold986/X _08628_/A2 _08618_/X _09977_/A sky130_fd_sc_hd__o211a_1
X_09599_ VGND VPWR VPWR VGND _14469_/D fanout70/X _09619_/S hold658/X sky130_fd_sc_hd__mux2_1
X_11630_ VGND VPWR VGND VPWR _11630_/X _12101_/A1 _11625_/X _11629_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
X_11561_ VPWR VGND VGND VPWR _11561_/A _11561_/Y _11561_/B sky130_fd_sc_hd__nand2_1
X_14080__1197 VPWR VGND VPWR VGND _15499_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
XFILLER_11_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10512_ VGND VPWR VGND VPWR _10512_/X _14946_/Q _10633_/A2 _10511_/X _10523_/A1 sky130_fd_sc_hd__o211a_1
X_11492_ VGND VPWR VPWR VGND _15081_/D _11491_/X _11492_/S _15081_/Q sky130_fd_sc_hd__mux2_1
X_14280_ hold535/A _14280_/CLK _14280_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10443_ VGND VPWR VPWR VGND _10443_/X hold765/A _10554_/S hold191/A sky130_fd_sc_hd__mux2_1
XFILLER_40_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10374_ VGND VPWR VGND VPWR _10374_/X _15006_/Q _10629_/A2 _10373_/X _10677_/S sky130_fd_sc_hd__o211a_1
X_12113_ VPWR VGND VGND VPWR _12113_/X hold202/A _12117_/B sky130_fd_sc_hd__or2_1
X_12944__61 VPWR VGND VPWR VGND _14187_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_12044_ VGND VPWR VGND VPWR _12044_/X hold995/A _12188_/A2 _11925_/S _12043_/X sky130_fd_sc_hd__o211a_1
XFILLER_78_777 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout790 VPWR VGND _09007_/A _08983_/A VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_65_427 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_1_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_19_811 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_clk clkload36/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_61_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_34_836 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_73_493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12877_ VGND VPWR VPWR VGND _15601_/D _07561_/X _12877_/S _07714_/A sky130_fd_sc_hd__mux2_1
X_15596_ _15596_/Q clkload55/A _15596_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11828_ VGND VPWR VPWR VGND _11828_/X hold969/A _11838_/S hold474/A sky130_fd_sc_hd__mux2_1
X_14616_ hold760/A _14616_/CLK _14616_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14547_ hold522/A _14547_/CLK _14547_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13487__604 VPWR VGND VPWR VGND _14762_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_11759_ VGND VPWR VPWR VGND _11759_/X _11756_/X _12098_/A _11755_/X sky130_fd_sc_hd__mux2_1
X_14478_ hold863/A _14478_/CLK _14478_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13528__645 VPWR VGND VPWR VGND _14808_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
XFILLER_66_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08970_ VGND VPWR VGND VPWR _15114_/D hold543/X _08985_/A2 _08969_/X _08943_/A sky130_fd_sc_hd__o211a_1
X_07921_ VPWR VGND VGND VPWR _07921_/A _07922_/B _07943_/A sky130_fd_sc_hd__nand2_1
X_07852_ VPWR VGND VPWR VGND clone18/X _15354_/Q _08495_/A2 _07852_/X _15143_/Q sky130_fd_sc_hd__a22o_1
Xinput1 VGND VPWR input1/X rst_n VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_56_438 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07783_ _08126_/B _07747_/X _07783_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_09522_ VPWR VGND VPWR VGND _09522_/Y _09549_/S sky130_fd_sc_hd__inv_2
XFILLER_37_641 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_clk clkload40/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_13080__197 VPWR VGND VPWR VGND _14323_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
XFILLER_80_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09453_ VPWR VGND VGND VPWR _09453_/X _09453_/A _09482_/S sky130_fd_sc_hd__or2_1
XFILLER_52_666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09384_ VGND VPWR VPWR VGND _14665_/D hold577/X _09411_/S clone133/X sky130_fd_sc_hd__mux2_1
X_08404_ VGND VPWR VPWR VGND _15373_/D _09548_/A1 _08411_/S hold486/X sky130_fd_sc_hd__mux2_1
XFILLER_40_839 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08335_ VGND VPWR VPWR VGND _15484_/D _09690_/A0 _08335_/S hold997/X sky130_fd_sc_hd__mux2_1
X_14201__919 _14201_/D _14201__919/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08266_ VGND VPWR VGND VPWR _08266_/X _08299_/A2 _15608_/Q _08255_/X _08265_/Y sky130_fd_sc_hd__a211o_2
X_08197_ VGND VPWR VPWR VGND _08197_/X _08193_/X _08197_/S _08195_/C sky130_fd_sc_hd__mux2_1
X_07217_ VGND VPWR _08223_/A _07368_/A _12845_/A VPWR VGND sky130_fd_sc_hd__xnor2_2
X_07148_ VPWR VGND VPWR VGND _08287_/A _07148_/A sky130_fd_sc_hd__inv_2
X_10090_ VPWR VGND VPWR VGND _10089_/X _10608_/A1 _10088_/X _10090_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_928 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_75_736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13321__438 VPWR VGND VPWR VGND _14596_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_39_clk clkload54/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12800_ VGND VPWR VPWR VGND _15557_/D _12799_/X _12798_/Y _12807_/A1 _12807_/B1 _15557_/Q
+ sky130_fd_sc_hd__a32o_1
XFILLER_47_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_43_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10992_ VGND VPWR VGND VPWR _10992_/X _10991_/X _10990_/X _11004_/A1 _11235_/C1 sky130_fd_sc_hd__a211o_1
X_12731_ VGND VPWR VPWR VGND _12732_/B _12730_/Y _12731_/S _12722_/Y sky130_fd_sc_hd__mux2_1
XFILLER_37_1019 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15450_ VGND VPWR VGND VPWR _15450_/Q _15450_/D clkload11/A sky130_fd_sc_hd__dfxtp_4
X_12662_ VGND VPWR VGND VPWR _12662_/X _12661_/X _12660_/X _12662_/A1 _12662_/C1 sky130_fd_sc_hd__a211o_1
X_11613_ VGND VPWR VPWR VGND _11617_/B hold427/A _12097_/S hold548/A sky130_fd_sc_hd__mux2_1
X_14401_ _14401_/Q clkload35/A _14401_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12593_ VGND VPWR VPWR VGND _12593_/X hold691/A _12599_/S _15058_/Q sky130_fd_sc_hd__mux2_1
X_13215__332 VPWR VGND VPWR VGND _14490_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_15381_ hold756/A _15381_/CLK _15381_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11544_ VPWR VGND VGND VPWR _11545_/B _15432_/D _11544_/B sky130_fd_sc_hd__nand2_1
X_14332_ hold682/A _14332_/CLK _14332_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14263_ hold771/A _14263_/CLK _14263_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11475_ VGND VPWR VPWR VGND _11475_/X _15077_/Q _11475_/S _15075_/Q sky130_fd_sc_hd__mux2_1
X_10426_ VGND VPWR VPWR VGND _10426_/X _10425_/X _10652_/S _10424_/X sky130_fd_sc_hd__mux2_1
X_14194_ _14194_/Q _14194_/CLK _14194_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10357_ VPWR VGND VPWR VGND _10356_/X _10608_/A1 _10355_/X _10357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_1304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10288_ VGND VPWR VPWR VGND _10288_/X _10287_/X _10288_/S _10286_/X sky130_fd_sc_hd__mux2_1
X_12027_ VPWR VGND VPWR VGND _12026_/X _12185_/A1 _12025_/X _12027_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_438 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_1286 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13903__1020 VPWR VGND VPWR VGND _15275_/CLK clkload13/A sky130_fd_sc_hd__inv_2
XFILLER_61_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15579_ _15579_/Q clkload31/A _15579_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08120_ VGND VPWR VGND VPWR _08120_/X _08182_/S _08116_/Y _08119_/X _08280_/B2 sky130_fd_sc_hd__o211a_1
X_08051_ VPWR VGND VPWR VGND _08051_/B _08051_/C _08051_/A _08051_/X sky130_fd_sc_hd__or3_1
X_13762__879 VPWR VGND VPWR VGND _15134_/CLK clkload19/A sky130_fd_sc_hd__inv_2
X_08953_ VPWR VGND _15120_/D _08953_/B _08955_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07904_ VGND VPWR VGND VPWR _07904_/X _10074_/A0 _07901_/X _07311_/B _07903_/Y sky130_fd_sc_hd__a211o_1
X_08884_ VPWR VGND VGND VPWR _08884_/X _15150_/Q _08926_/B sky130_fd_sc_hd__or2_1
XFILLER_56_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07835_ VGND VPWR VGND VPWR _08059_/B _08145_/A _15552_/Q _15553_/Q _15554_/Q sky130_fd_sc_hd__and4_2
X_07766_ VPWR VGND VPWR VGND _07769_/C _07769_/B _07769_/A _07766_/Y sky130_fd_sc_hd__a21oi_1
X_13656__773 VPWR VGND VPWR VGND _14996_/CLK clkload38/A sky130_fd_sc_hd__inv_2
XFILLER_53_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09505_ VGND VPWR VPWR VGND _14554_/D fanout29/X _09513_/S hold745/X sky130_fd_sc_hd__mux2_1
X_07697_ VPWR VGND VPWR VGND _07695_/X _07694_/A _07414_/Y _07697_/X _08225_/C1 sky130_fd_sc_hd__a22o_1
X_09436_ VGND VPWR VPWR VGND _14616_/D fanout19/X _09441_/S hold760/X sky130_fd_sc_hd__mux2_1
XFILLER_52_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09367_ VGND VPWR VPWR VGND _14679_/D hold504/X _09379_/S fanout17/X sky130_fd_sc_hd__mux2_1
X_08318_ VGND VPWR VPWR VGND _15501_/D fanout44/X _08318_/S hold963/X sky130_fd_sc_hd__mux2_1
X_09298_ VGND VPWR VPWR VGND _14743_/D fanout16/X _09310_/S hold659/X sky130_fd_sc_hd__mux2_1
XANTENNA_50 _10505_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_72 _09790_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_83 _08190_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08249_ VPWR VGND VPWR VGND _08245_/X _15609_/Q _08249_/A2 _08250_/A _08249_/B2 sky130_fd_sc_hd__a22o_1
XANTENNA_61 _09414_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_94 _14407_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11260_ VGND VPWR VPWR VGND _11260_/X _15194_/Q _11261_/B _15062_/Q sky130_fd_sc_hd__mux2_1
X_12914__31 VPWR VGND VPWR VGND _14157_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
XFILLER_49_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10211_ VPWR VGND VGND VPWR _11210_/A _10211_/B _10211_/Y sky130_fd_sc_hd__nor2_1
X_11191_ VPWR VGND VPWR VGND _11190_/X _11173_/A _12713_/B1 _11191_/X sky130_fd_sc_hd__a21o_1
X_10142_ VGND VPWR VPWR VGND _10142_/X hold983/A _10604_/S hold702/A sky130_fd_sc_hd__mux2_1
X_10073_ VPWR VGND VPWR VGND _10071_/C _10071_/B _11535_/C _10073_/Y sky130_fd_sc_hd__a21oi_1
X_14950_ hold828/A _14950_/CLK _14950_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14881_ _14881_/Q _14881_/CLK _14881_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1321 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15502_ _15502_/Q _15502_/CLK _15502_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_43_452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12714_ VPWR VGND VGND VPWR _12695_/Y _12713_/X _12751_/A2 _15475_/Q _15475_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
X_10975_ VPWR VGND VGND VPWR _10975_/X _10995_/S _10975_/B sky130_fd_sc_hd__or2_1
XFILLER_43_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15433_ _15433_/Q clkload47/A _15433_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12645_ VPWR VGND VGND VPWR _12645_/X _12655_/S _12645_/B sky130_fd_sc_hd__or2_1
X_15364_ hold150/A _15364_/CLK _15364_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12576_ VGND VPWR VPWR VGND _12576_/X _14278_/Q _12594_/B _14310_/Q sky130_fd_sc_hd__mux2_1
XFILLER_62_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11527_ VGND VPWR VPWR VGND _11527_/X _11526_/X _11530_/S _15473_/Q sky130_fd_sc_hd__mux2_1
X_14315_ hold602/A _14315_/CLK _14315_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15295_ _15295_/Q _15295_/CLK _15295_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14246_ _14246_/Q _14246_/CLK _14246_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11458_ VGND VPWR VPWR VGND _11458_/X _11457_/X _11458_/S _15450_/Q sky130_fd_sc_hd__mux2_1
Xhold309 hold309/X hold309/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11389_ VPWR VGND VGND VPWR _11389_/X _14818_/Q _11392_/B sky130_fd_sc_hd__or2_1
X_10409_ VGND VPWR VPWR VGND _10409_/X hold399/A _10702_/S hold616/A sky130_fd_sc_hd__mux2_1
X_14177_ hold628/A _14177_/CLK _14177_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13599__716 VPWR VGND VPWR VGND _14939_/CLK clkload35/A sky130_fd_sc_hd__inv_2
XFILLER_78_371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1009 hold1009/X _15272_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13343__460 VPWR VGND VPWR VGND _14618_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_6_1326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_1189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07620_ VGND VPWR _07620_/B _07620_/Y _07625_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07551_ VPWR VGND VGND VPWR _07551_/X _07551_/A _07551_/B sky130_fd_sc_hd__or2_1
XFILLER_35_920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07482_ VPWR VGND VGND VPWR _07483_/B _15447_/Q _07482_/B sky130_fd_sc_hd__or2_1
XFILLER_50_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09221_ VGND VPWR VPWR VGND _14872_/D hold781/X _09231_/S fanout10/X sky130_fd_sc_hd__mux2_1
X_09152_ VGND VPWR VPWR VGND _14946_/D _08091_/X _09163_/S hold1084/X sky130_fd_sc_hd__mux2_1
X_08103_ VGND VPWR VGND VPWR _08103_/X _08277_/S _10063_/B _08101_/Y _08280_/B2 sky130_fd_sc_hd__o211a_1
X_09083_ VGND VPWR VPWR VGND _15010_/D hold1135/X _09094_/S fanout13/X sky130_fd_sc_hd__mux2_1
X_08034_ VPWR VGND VPWR VGND _08034_/B1 _15345_/Q _08253_/A2 _08034_/X _15150_/Q sky130_fd_sc_hd__a22o_1
Xhold821 hold821/X hold821/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold810 hold810/X hold810/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 hold854/X hold854/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 hold832/X hold832/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 hold843/X hold843/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 hold865/X hold865/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 hold887/X hold887/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 hold876/X hold876/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 hold898/X hold898/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ VPWR VGND _09989_/C _09986_/B _15609_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_08936_ VPWR VGND VGND VPWR _09873_/A _15479_/Q _09869_/A _08936_/X sky130_fd_sc_hd__o21a_1
X_08867_ VGND VPWR VGND VPWR _15159_/D hold1181/X _08893_/A2 _08866_/X _09024_/A sky130_fd_sc_hd__o211a_1
X_07818_ VGND VPWR _07878_/B _07859_/A _07856_/A _07855_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
X_08798_ VGND VPWR VPWR VGND _15211_/D fanout31/X _08814_/S hold230/X sky130_fd_sc_hd__mux2_1
X_13392__509 VPWR VGND VPWR VGND _14667_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_07749_ VPWR VGND VPWR VGND _07751_/C _15598_/Q _15551_/Q _07750_/B sky130_fd_sc_hd__a21o_1
XFILLER_26_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14207__925 _14207_/D _14207__925/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_10760_ VGND VPWR VPWR VGND _10760_/X hold867/A _10835_/B hold508/A sky130_fd_sc_hd__mux2_1
X_10691_ VGND VPWR VPWR VGND _10691_/X hold998/A _10702_/S hold536/A sky130_fd_sc_hd__mux2_1
X_09419_ VGND VPWR VPWR VGND _14633_/D fanout84/X _09446_/S hold500/X sky130_fd_sc_hd__mux2_1
X_12430_ VGND VPWR VPWR VGND _12430_/X hold716/A _12651_/S hold251/A sky130_fd_sc_hd__mux2_1
X_12361_ VGND VPWR VPWR VGND _12361_/X hold823/A _12599_/S hold697/A sky130_fd_sc_hd__mux2_1
X_13286__403 VPWR VGND VPWR VGND _14561_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_11312_ VPWR VGND VGND VPWR _11421_/C _11313_/C _11421_/B sky130_fd_sc_hd__nor2_2
X_13979__1096 VPWR VGND VPWR VGND _15351_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_12292_ VPWR VGND VGND VPWR _12292_/X hold585/A _12701_/S sky130_fd_sc_hd__or2_1
X_15080_ _15080_/Q clkload37/A _15080_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_4_323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11243_ VGND VPWR VGND VPWR _11243_/X _11252_/C1 _11239_/X _11242_/X _11254_/C1 sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_26_Left_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13327__444 VPWR VGND VPWR VGND _14602_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_80_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11174_ VGND VPWR VPWR VGND _11174_/X _14440_/Q _11175_/S _14696_/Q sky130_fd_sc_hd__mux2_1
XFILLER_48_511 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10125_ VGND VPWR VGND VPWR _10125_/X _10347_/A1 _10121_/X _10124_/X _10622_/C1 sky130_fd_sc_hd__o211a_1
X_14933_ _14933_/Q clkload30/A _14933_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_62_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10056_ VPWR VGND VGND VPWR _10056_/A _11340_/A _10056_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_72 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_23_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14864_ hold927/A _14864_/CLK _14864_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_35_Left_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14795_ _14795_/Q _14795_/CLK _14795_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10958_ VGND VPWR VGND VPWR _10958_/X _10957_/X _10956_/X _11170_/S _11180_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_16_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15416_ hold452/A _15416_/CLK _15416_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10889_ VGND VPWR VGND VPWR _10889_/X _10890_/A _10885_/X _10888_/X _12868_/A1 sky130_fd_sc_hd__o211a_1
X_12628_ VGND VPWR VGND VPWR _12628_/X _12627_/X _12626_/X _12624_/S _12739_/C1 sky130_fd_sc_hd__a211o_1
X_15347_ _15347_/Q _15347_/CLK _15347_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12559_ VGND VPWR VGND VPWR _12559_/X _12556_/X _12558_/X _12674_/A1 _12740_/A1 sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_44_Left_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15278_ _15278_/Q _15278_/CLK _15278_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14229_ hold189/A _14229_/CLK _14229_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout608 VGND VPWR _08377_/Y _08408_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout619 _09867_/S _09865_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_28_1349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09770_ VGND VPWR VPWR VGND _14279_/D _09792_/S fanout76/X hold1214/X sky130_fd_sc_hd__mux2_4
X_08721_ VGND VPWR VGND VPWR _15273_/D hold840/X _08721_/A2 _08720_/X _11294_/A sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_53_Left_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08652_ VPWR VGND VPWR VGND _15294_/Q _08714_/A2 _08652_/X _08711_/B1 _08651_/X _08722_/C1
+ sky130_fd_sc_hd__a221o_1
X_07603_ VPWR VGND VPWR VGND _15135_/Q clone20/X _15362_/Q _08253_/A2 _07603_/X sky130_fd_sc_hd__a22o_2
X_08583_ VGND VPWR VGND VPWR _08583_/X _08617_/A _08615_/B1 hold989/X _08582_/Y sky130_fd_sc_hd__a211o_1
X_13120__237 VPWR VGND VPWR VGND _14363_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_39_1412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07534_ VPWR VGND VGND VPWR _07534_/A _07534_/B _07534_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07465_ VGND VPWR VPWR VGND _07467_/B _09240_/A _07469_/S _15594_/Q sky130_fd_sc_hd__mux2_1
X_09204_ VGND VPWR VPWR VGND _14889_/D _09228_/S hold1212/X fanout73/X sky130_fd_sc_hd__mux2_4
X_13768__885 VPWR VGND VPWR VGND _15140_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_07396_ VPWR VGND VPWR VGND _07395_/X _07820_/A _07391_/X _07397_/C sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_62_Left_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09135_ VGND VPWR VPWR VGND _14963_/D _09157_/S clone146/X hold1269/X sky130_fd_sc_hd__mux2_4
X_13014__131 VPWR VGND VPWR VGND _14257_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_09066_ VGND VPWR VPWR VGND _15027_/D hold1088/X _09090_/S fanout77/X sky130_fd_sc_hd__mux2_1
X_08017_ VGND VPWR VPWR VGND _08017_/X _08016_/X _08195_/A _07603_/X sky130_fd_sc_hd__mux2_1
Xhold651 hold651/X hold651/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_838 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold640 hold640/X hold640/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 hold662/X hold662/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 hold684/X hold684/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 hold695/X hold695/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 hold673/X hold673/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09968_ VPWR VGND VPWR VGND _14801_/Q _09966_/X _14801_/D _09967_/Y _10060_/A _11340_/A
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_71_Left_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08919_ VGND VPWR VGND VPWR _15133_/D hold1186/X _08919_/A2 _08918_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
X_09899_ VGND VPWR _08859_/C hold714/A _09900_/B _14144_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold1340 hold1340/X _15352_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1351 hold1351/X _14998_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11930_ VGND VPWR VGND VPWR _11930_/X _11927_/X _11929_/X _12156_/A1 _12202_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_79_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1373 hold1373/X _15139_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 _10042_/A _15633_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 hold1395/X _15084_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _09593_/A _14474_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11861_ VPWR VGND _11861_/X _11860_/X _11856_/X _12102_/S _11852_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11792_ VGND VPWR VPWR VGND _11792_/X hold805/A _12589_/S hold279/A sky130_fd_sc_hd__mux2_1
X_10812_ VGND VPWR VPWR VGND _10816_/B hold881/A _11223_/S hold209/A sky130_fd_sc_hd__mux2_1
X_14580_ hold330/A _14580_/CLK _14580_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10743_ VPWR VGND VGND VPWR _10743_/X hold622/A _10743_/B sky130_fd_sc_hd__or2_1
XFILLER_43_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15201_ hold243/A _15201_/CLK _15201_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10674_ VPWR VGND VGND VPWR _10655_/Y _10673_/X _10562_/B _14394_/Q _14394_/D _12159_/C1
+ sky130_fd_sc_hd__o221a_1
X_12413_ VPWR VGND VGND VPWR _12413_/X hold589/A _12726_/S sky130_fd_sc_hd__or2_1
X_12344_ VPWR VGND VGND VPWR _12325_/Y _12343_/X _12269_/B _15465_/Q _15465_/D _11341_/A
+ sky130_fd_sc_hd__o221a_1
X_15132_ _15132_/Q _15132_/CLK _15132_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15063_ _15063_/Q _15063_/CLK _15063_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12275_ VPWR VGND VGND VPWR _12275_/X _12698_/S _12275_/B sky130_fd_sc_hd__or2_1
X_13561__678 VPWR VGND VPWR VGND _14892_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_11226_ VGND VPWR VGND VPWR _11226_/X _11223_/X _11225_/X _10816_/A _11263_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_4_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11157_ VGND VPWR VPWR VGND _11157_/X _14504_/Q _11167_/S _14184_/Q sky130_fd_sc_hd__mux2_1
X_10108_ VGND VPWR VGND VPWR _10108_/X _10608_/A1 _10103_/X _10107_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
X_11088_ VGND VPWR VGND VPWR _11088_/X _11087_/X _11086_/X _11092_/S _11217_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_27_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10039_ VPWR VGND VPWR VGND _10038_/C _15631_/Q hold1308/X _10040_/B sky130_fd_sc_hd__a21oi_1
X_14916_ _14916_/Q _14916_/CLK _14916_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14847_ _14847_/Q clkload20/A _14847_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13455__572 VPWR VGND VPWR VGND _14730_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_14778_ hold879/A _14778_/CLK _14778_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07250_ VPWR VGND VGND VPWR _14391_/Q _07230_/S _07265_/B1 _07252_/B sky130_fd_sc_hd__o21a_1
X_07181_ VPWR VGND VPWR VGND _07181_/Y _07972_/A sky130_fd_sc_hd__inv_2
XFILLER_69_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13802__919 VPWR VGND VPWR VGND _15174_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_14049__1166 VPWR VGND VPWR VGND _15421_/CLK clkload42/A sky130_fd_sc_hd__inv_2
Xfanout405 VGND VPWR fanout405/A _10846_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout438 VGND VPWR _11096_/C1 _11263_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout427 VPWR VGND _10634_/C1 _10505_/A1 VPWR VGND sky130_fd_sc_hd__buf_4
X_09822_ VGND VPWR VPWR VGND _14230_/D fanout12/X _09833_/S hold360/X sky130_fd_sc_hd__mux2_1
Xfanout416 VGND VPWR _12868_/A1 _10918_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout449 VPWR VGND _10626_/C1 _10737_/C1 VPWR VGND sky130_fd_sc_hd__buf_4
X_09753_ VGND VPWR VPWR VGND _14293_/D fanout8/X _09763_/S hold176/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08704_ VGND VPWR VGND VPWR _15280_/D hold1213/X _08704_/A2 _08703_/X _12159_/C1
+ sky130_fd_sc_hd__o211a_1
X_09684_ VGND VPWR VPWR VGND _14356_/D hold981/X _09684_/S fanout6/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_867 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08635_ VPWR VGND VGND VPWR _08635_/X _14393_/Q _08640_/B sky130_fd_sc_hd__or2_1
X_13978__1095 VPWR VGND VPWR VGND _15350_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_08566_ VPWR VGND _08566_/X _08566_/B _08566_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07517_ VGND VPWR _15465_/Q _07519_/B _07539_/C _15466_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xfanout12 VGND VPWR fanout13/X fanout12/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_08497_ VPWR VGND VPWR VGND _14135_/Q hold539/A _14134_/Q _14136_/Q _08500_/C sky130_fd_sc_hd__or4_1
Xfanout45 VGND VPWR _07910_/X fanout45/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout34 VGND VPWR _07994_/X fanout34/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout56 VPWR VGND VGND VPWR clone55/A fanout56/X sky130_fd_sc_hd__buf_8
Xfanout23 VPWR VGND VGND VPWR fanout24/X fanout23/X sky130_fd_sc_hd__buf_8
X_07448_ VPWR VGND _07450_/A _11535_/A _15455_/Q VPWR VGND sky130_fd_sc_hd__and2_1
Xfanout89 VPWR VGND VGND VPWR fanout90/X fanout89/X sky130_fd_sc_hd__buf_8
Xfanout67 VGND VPWR _07688_/X fanout67/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout78 VPWR VGND fanout78/X fanout79/X VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_52_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07379_ VPWR VGND VGND VPWR _07254_/Y _07357_/Y _07356_/Y _08081_/A _08081_/B _07379_/X
+ sky130_fd_sc_hd__a311o_2
X_09118_ VGND VPWR VPWR VGND _14977_/D hold391/X _09128_/S fanout10/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10390_ VGND VPWR VPWR VGND _10390_/X hold569/A _10390_/S hold615/A sky130_fd_sc_hd__mux2_1
X_09049_ VGND VPWR VPWR VGND _15041_/D hold788/X _09059_/S fanout9/A sky130_fd_sc_hd__mux2_1
XFILLER_78_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold470 hold470/X hold470/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12060_ VGND VPWR VPWR VGND _12060_/X hold744/A _12219_/S hold444/A sky130_fd_sc_hd__mux2_1
XFILLER_1_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold481 hold481/X hold481/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 hold492/X hold492/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ VGND VPWR VPWR VGND _11011_/X hold740/A _11165_/S hold467/A sky130_fd_sc_hd__mux2_1
X_13398__515 VPWR VGND VPWR VGND _14673_/CLK clkload54/A sky130_fd_sc_hd__inv_2
XFILLER_65_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1170 hold1170/X _14305_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1192 _07123_/A _15477_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_642 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1181 hold1181/X _15158_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14701_ hold401/A _14701_/CLK _14701_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13439__556 VPWR VGND VPWR VGND _14714_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_11913_ VPWR VGND VGND VPWR _11913_/X _12069_/S _11913_/B sky130_fd_sc_hd__or2_1
XFILLER_79_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11844_ VPWR VGND VGND VPWR _12103_/A _11844_/B _11844_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14632_ _14632_/Q _14632_/CLK _14632_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11775_ VGND VPWR VGND VPWR _11775_/X hold856/A _12188_/A2 _12008_/A1 _11774_/X sky130_fd_sc_hd__o211a_1
X_14563_ hold516/A _14563_/CLK _14563_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14494_ _14494_/Q _14494_/CLK _14494_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10726_ VGND VPWR VPWR VGND _10726_/X _10723_/X _10732_/S _10722_/X sky130_fd_sc_hd__mux2_1
X_10657_ VGND VPWR VGND VPWR _10657_/X _14877_/Q _10744_/A2 _10656_/X _10652_/S sky130_fd_sc_hd__o211a_1
Xclkload26 VGND VPWR VGND VPWR clkload26/A clkload26/Y sky130_fd_sc_hd__clkinv_8
Xclkload15 clkload15/Y clkload15/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload48 clkload48/Y clkload48/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload37 clkload37/Y clkload37/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
X_10588_ VGND VPWR VPWR VGND _10588_/X _10587_/X _10588_/S _10586_/X sky130_fd_sc_hd__mux2_1
X_15115_ hold888/A _15115_/CLK _15115_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12327_ VGND VPWR VPWR VGND _12327_/X hold880/A _12339_/B hold652/A sky130_fd_sc_hd__mux2_1
X_12258_ VGND VPWR VPWR VGND _12262_/B hold726/A _12339_/B hold432/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15046_ hold660/A _15046_/CLK _15046_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11209_ VGND VPWR VPWR VGND _11210_/B _11208_/Y _11209_/S _11200_/Y sky130_fd_sc_hd__mux2_1
X_12189_ VGND VPWR VGND VPWR _12189_/X _12186_/X _12188_/X _11894_/S _12189_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_49_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08420_ VPWR VGND VPWR VGND _08418_/X hold150/X _08419_/Y _15364_/D sky130_fd_sc_hd__a21oi_1
X_13191__308 VPWR VGND VPWR VGND _14466_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_08351_ VGND VPWR VPWR VGND _15422_/D hold711/X _08372_/S fanout62/X sky130_fd_sc_hd__mux2_1
X_08282_ VGND VPWR VPWR VGND _08282_/X _08273_/B _08273_/A _07810_/A _12833_/A _14153_/Q
+ sky130_fd_sc_hd__a32o_1
X_07302_ VPWR VGND VGND VPWR _07813_/A _07311_/A _07817_/A sky130_fd_sc_hd__nor2_1
X_07233_ VPWR VGND VPWR VGND _10061_/A _08257_/B _07221_/X _08239_/A sky130_fd_sc_hd__a21o_1
Xclkload9 VGND VPWR VPWR VGND clkload9/A clkload9/Y sky130_fd_sc_hd__clkinvlp_4
X_13232__349 VPWR VGND VPWR VGND _14507_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_07164_ VPWR VGND VGND VPWR _14406_/Q _07301_/A2 _07301_/B1 _07166_/B sky130_fd_sc_hd__o21a_1
X_07095_ VPWR VGND VPWR VGND _07368_/A _15449_/Q sky130_fd_sc_hd__inv_2
X_13085__202 VPWR VGND VPWR VGND _14328_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
Xfanout213 VGND VPWR fanout217/X _12748_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout202 VGND VPWR _12226_/A1 _11894_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout246 VGND VPWR _12666_/A1 _12656_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout235 VGND VPWR _12008_/C1 _12101_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout224 VPWR VGND _12226_/C1 fanout234/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout257 VPWR VGND _12176_/S _12139_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_07997_ VPWR VGND VGND VPWR _07570_/X _07421_/Y _12080_/A2 _07421_/A _08014_/A _07996_/X
+ sky130_fd_sc_hd__o221a_1
Xfanout268 VPWR VGND _12732_/A _07912_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout279 VGND VPWR fanout282/X _11184_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09805_ VGND VPWR VPWR VGND _14247_/D _09827_/S fanout76/X hold1180/X sky130_fd_sc_hd__mux2_4
X_13126__243 VPWR VGND VPWR VGND _14369_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_09736_ VGND VPWR VPWR VGND _14310_/D _09760_/S clone47/A hold1133/X sky130_fd_sc_hd__mux2_4
XFILLER_55_631 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09667_ VGND VPWR VPWR VGND _14373_/D hold783/X _09687_/S fanout69/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08618_ VGND VPWR VGND VPWR _08618_/X _08617_/A _08627_/C1 hold1079/X _08617_/Y sky130_fd_sc_hd__a211o_1
X_09598_ VGND VPWR VPWR VGND _14470_/D _09619_/S clone47/A hold1266/X sky130_fd_sc_hd__mux2_4
X_08549_ VGND VPWR _08548_/C _08548_/A _08549_/Y _08548_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_39_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11560_ VPWR VGND VPWR VGND _11559_/Y _11561_/B _11341_/Y _15440_/D sky130_fd_sc_hd__a21oi_1
X_13783__900 VPWR VGND VPWR VGND _15155_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_10511_ VPWR VGND VGND VPWR _10511_/X hold322/A _10516_/S sky130_fd_sc_hd__or2_1
X_11491_ VGND VPWR VPWR VGND _11491_/X _11490_/X _11491_/S _15461_/Q sky130_fd_sc_hd__mux2_1
X_13824__941 VPWR VGND VPWR VGND _15196_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_10442_ VGND VPWR VPWR VGND _10446_/B hold750/A _10554_/S hold158/A sky130_fd_sc_hd__mux2_1
X_10373_ VPWR VGND VGND VPWR _10373_/X hold524/A _10696_/S sky130_fd_sc_hd__or2_1
X_12112_ VGND VPWR VPWR VGND _12112_/X hold733/A _12112_/S hold300/A sky130_fd_sc_hd__mux2_1
X_12043_ VPWR VGND VGND VPWR _12043_/X hold899/A _12043_/B sky130_fd_sc_hd__or2_1
Xfanout791 VGND VPWR _15478_/Q _08983_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout780 VPWR VGND _07301_/B1 _07265_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_37_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_61_634 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12876_ VGND VPWR VPWR VGND _15600_/D _07603_/X _14802_/D hold1272/X sky130_fd_sc_hd__mux2_1
XFILLER_45_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15595_ _15595_/Q clkload45/A _15595_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11827_ VGND VPWR VPWR VGND _11831_/B hold462/A _11838_/S hold350/A sky130_fd_sc_hd__mux2_1
X_14615_ hold547/A _14615_/CLK _14615_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14048__1165 VPWR VGND VPWR VGND _15420_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_14546_ hold665/A _14546_/CLK _14546_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11758_ VGND VPWR VGND VPWR _11758_/X _12099_/A1 _11754_/X _11757_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
X_10709_ VPWR VGND VPWR VGND _10709_/X _10507_/A _10682_/X _10690_/X _10708_/X _10707_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_18_1167 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14477_ _14477_/Q _14477_/CLK _14477_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11689_ VGND VPWR VPWR VGND _11689_/X _14190_/Q _12479_/S hold190/A sky130_fd_sc_hd__mux2_1
X_13567__684 VPWR VGND VPWR VGND _14898_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_13977__1094 VPWR VGND VPWR VGND _15349_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_07920_ VGND VPWR _07942_/C _07945_/A _07943_/A _07942_/B VPWR VGND sky130_fd_sc_hd__o21ai_1
X_15029_ _15029_/Q _15029_/CLK _15029_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07851_ VGND VPWR VGND VPWR _15354_/Q _08495_/A2 _15143_/Q _07851_/Y _07873_/B1 sky130_fd_sc_hd__a22oi_4
Xinput2 VGND VPWR input2/X ui_in[0] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_12890__7 VPWR VGND VPWR VGND _14132_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_07782_ VPWR VGND VPWR VGND _07751_/C _15599_/Q _15552_/Q _07783_/B sky130_fd_sc_hd__a21o_1
XFILLER_42_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09521_ VPWR VGND _09521_/A _09521_/X _09834_/A VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_37_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09452_ VPWR VGND VPWR VGND _09452_/Y _09482_/S sky130_fd_sc_hd__inv_2
XFILLER_25_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_678 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08403_ VGND VPWR VPWR VGND _15374_/D _09547_/A1 _08409_/S hold680/X sky130_fd_sc_hd__mux2_1
X_09383_ _14666_/D fanout94/X fanout90/X _09411_/S _09382_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08334_ VGND VPWR VPWR VGND _15485_/D _09655_/A0 _08335_/S hold1050/X sky130_fd_sc_hd__mux2_1
X_13808__925 VPWR VGND VPWR VGND _15180_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_08265_ VGND VPWR VGND VPWR _08147_/A _08265_/Y _08220_/A _15545_/Q _08256_/X _08264_/Y
+ sky130_fd_sc_hd__o221ai_4
X_08196_ VPWR VGND VGND VPWR _08193_/X _08194_/Y _08035_/X _08194_/B _08196_/X _08195_/X
+ sky130_fd_sc_hd__o221a_1
X_07216_ VPWR VGND _07216_/X _12845_/A _15449_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07147_ VPWR VGND VGND VPWR _07148_/A _15476_/Q _07149_/B sky130_fd_sc_hd__or2_1
XFILLER_10_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13360__477 VPWR VGND VPWR VGND _14635_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XFILLER_55_461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09719_ VGND VPWR VPWR VGND _14324_/D fanout6/X _09721_/S hold773/X sky130_fd_sc_hd__mux2_1
X_10991_ VGND VPWR VPWR VGND _10991_/X hold729/A _11241_/S hold382/A sky130_fd_sc_hd__mux2_1
X_12730_ VPWR VGND VPWR VGND _12729_/X _12740_/A1 _12728_/X _12730_/Y sky130_fd_sc_hd__a21oi_1
X_12661_ VGND VPWR VPWR VGND _12661_/X hold813/A _12661_/S hold424/A sky130_fd_sc_hd__mux2_1
X_14400_ _14400_/Q clkload44/A _14400_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11612_ VPWR VGND VPWR VGND _11611_/X _12008_/C1 _11610_/X _11612_/Y sky130_fd_sc_hd__a21oi_1
X_12592_ VGND VPWR VGND VPWR _12592_/X _12744_/C1 _12591_/X _12588_/X _12864_/A1 sky130_fd_sc_hd__o211a_1
X_15380_ hold733/A _15380_/CLK _15380_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13254__371 VPWR VGND VPWR VGND _14529_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_11543_ VPWR VGND VPWR VGND _11269_/B hold1144/X _11542_/A _11544_/B sky130_fd_sc_hd__a21oi_1
X_14331_ hold938/A _14331_/CLK _14331_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11474_ VGND VPWR VPWR VGND _15075_/D _11473_/X _11477_/S _15075_/Q sky130_fd_sc_hd__mux2_1
X_14262_ hold459/A _14262_/CLK _14262_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14193_ _14193_/Q _14193_/CLK _14193_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10425_ VGND VPWR VPWR VGND _10425_/X hold538/A _10720_/S hold312/A sky130_fd_sc_hd__mux2_1
X_10356_ VGND VPWR VPWR VGND _10356_/X _10353_/X _10615_/S _10352_/X sky130_fd_sc_hd__mux2_1
X_13601__718 VPWR VGND VPWR VGND _14941_/CLK clkload55/A sky130_fd_sc_hd__inv_2
XFILLER_3_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10287_ VGND VPWR VPWR VGND _10287_/X hold779/A _10664_/S hold494/A sky130_fd_sc_hd__mux2_1
X_12026_ VGND VPWR VPWR VGND _12026_/X _12023_/X _12180_/S _12022_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_46_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_59_1256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_995 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12859_ VGND VPWR VPWR VGND _15583_/D _08034_/X _12860_/S _07331_/A sky130_fd_sc_hd__mux2_1
X_15578_ _15578_/Q clkload32/A _15578_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14529_ hold168/A _14529_/CLK _14529_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08050_ VPWR VGND VPWR VGND _08049_/Y _08046_/X _10059_/A _08051_/C sky130_fd_sc_hd__a21oi_1
X_08952_ VPWR VGND VPWR VGND _08969_/A _15119_/Q _08933_/A _08953_/B _15120_/Q sky130_fd_sc_hd__a22o_1
X_08883_ VGND VPWR VGND VPWR _15151_/D hold1161/X _08919_/A2 _08882_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
X_07903_ VGND VPWR _10075_/A _07902_/X _07903_/Y _07899_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_57_737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07834_ VPWR VGND VGND VPWR _15552_/Q _08099_/B _08145_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07765_ VPWR VGND VGND VPWR _15592_/Q _07769_/C _07765_/B sky130_fd_sc_hd__nand2_1
X_13197__314 VPWR VGND VPWR VGND _14472_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
XFILLER_77_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09504_ VGND VPWR VPWR VGND _14555_/D fanout32/X _09520_/S hold613/X sky130_fd_sc_hd__mux2_1
X_07696_ VGND VPWR VGND VPWR _07668_/B _07316_/B _07972_/B _07696_/X _07316_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09435_ VGND VPWR VPWR VGND _14617_/D fanout23/X _09449_/S hold521/X sky130_fd_sc_hd__mux2_1
X_13238__355 VPWR VGND VPWR VGND _14513_/CLK clkload55/A sky130_fd_sc_hd__inv_2
XFILLER_52_486 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09366_ VGND VPWR VPWR VGND _14680_/D hold799/X _09377_/S fanout20/X sky130_fd_sc_hd__mux2_1
XANTENNA_40 _12213_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08317_ VGND VPWR VPWR VGND _08332_/S fanout49/X hold1196/X _15502_/D sky130_fd_sc_hd__mux2_2
X_09297_ VGND VPWR VPWR VGND _14744_/D fanout19/X _09302_/S hold444/X sky130_fd_sc_hd__mux2_1
XANTENNA_84 _08377_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08248_ VPWR VGND VGND VPWR _08147_/A _08246_/Y _08220_/A _08247_/X _08248_/X sky130_fd_sc_hd__o22a_1
XANTENNA_62 _09377_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_73 _09790_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_51 _10505_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_95 _14407_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08179_ VGND VPWR VPWR VGND _08180_/A _12766_/B _08179_/B sky130_fd_sc_hd__xor2_1
X_10210_ VGND VPWR VPWR VGND _10211_/B _10209_/Y _10987_/S _10201_/Y sky130_fd_sc_hd__mux2_1
X_11190_ VPWR VGND _11190_/X _11189_/X _11185_/X _11209_/S _11181_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14047__1164 VPWR VGND VPWR VGND _15419_/CLK clkload47/A sky130_fd_sc_hd__inv_2
XFILLER_0_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10141_ VGND VPWR VGND VPWR _10141_/X _10140_/X _10139_/X _10347_/A1 _10614_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_43_1002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10072_ VPWR VGND VGND VPWR _10072_/A _10072_/Y _10072_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_75_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14880_ hold868/A _14880_/CLK _14880_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_75_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_56_770 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10974_ VGND VPWR VPWR VGND _10974_/X hold516/A _10994_/S hold269/A sky130_fd_sc_hd__mux2_1
X_13976__1093 VPWR VGND VPWR VGND _15348_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_15501_ hold963/A _15501_/CLK _15501_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12713_ VPWR VGND VPWR VGND _12712_/X _12732_/A _12713_/B1 _12713_/X sky130_fd_sc_hd__a21o_1
X_15432_ _15432_/Q clkload47/A _15432_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12644_ VGND VPWR VPWR VGND _12644_/X hold580/A _12651_/S hold403/A sky130_fd_sc_hd__mux2_1
X_12575_ VGND VPWR VPWR VGND _12579_/B _14795_/Q _12577_/S _14246_/Q sky130_fd_sc_hd__mux2_1
X_15363_ _15363_/Q _15363_/CLK _15363_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11526_ VGND VPWR VPWR VGND _11526_/X _15094_/Q _11529_/S _15092_/Q sky130_fd_sc_hd__mux2_1
X_14314_ _14314_/Q _14314_/CLK _14314_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15294_ _15294_/Q _15294_/CLK _15294_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11457_ VGND VPWR VPWR VGND _11457_/X _15071_/Q _11490_/S _15069_/Q sky130_fd_sc_hd__mux2_1
X_14245_ hold283/A _14245_/CLK _14245_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13031__148 VPWR VGND VPWR VGND _14274_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_14176_ hold405/A _14176_/CLK _14176_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11388_ VGND VPWR VPWR VGND _14849_/D _11387_/X _11388_/S hold1299/X sky130_fd_sc_hd__mux2_1
X_10408_ VGND VPWR VGND VPWR _10408_/X _10405_/X _10407_/X _10705_/A _10704_/C1 sky130_fd_sc_hd__a211o_1
X_10339_ VPWR VGND VPWR VGND _10339_/X _11173_/A _10312_/X _10320_/X _10338_/X _10337_/X
+ sky130_fd_sc_hd__o32a_1
X_13679__796 VPWR VGND VPWR VGND _15019_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_12009_ VPWR VGND _12009_/X _12008_/X _12004_/X _12102_/S _12000_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_38_214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07550_ VPWR VGND _07560_/C _07556_/B _08956_/B VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_47_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_59_1042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07481_ VPWR VGND VGND VPWR _07479_/Y _07573_/A _07476_/Y _07580_/A sky130_fd_sc_hd__o21a_1
XFILLER_35_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09220_ VGND VPWR VPWR VGND _14873_/D hold994/X _09231_/S fanout13/X sky130_fd_sc_hd__mux2_1
X_09151_ VGND VPWR VPWR VGND _14947_/D fanout15/X _09163_/S hold637/X sky130_fd_sc_hd__mux2_1
X_08102_ VGND VPWR _08102_/B _10063_/B _08102_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_09082_ VGND VPWR VPWR VGND _15011_/D hold995/X _09094_/S _08070_/X sky130_fd_sc_hd__mux2_1
X_08033_ VGND VPWR VPWR VGND _15527_/D fanout25/X _08300_/S hold300/X sky130_fd_sc_hd__mux2_1
Xhold811 hold811/X hold811/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold800 hold800/X hold800/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 hold855/X hold855/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 hold844/X hold844/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 hold822/X hold822/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 hold833/X hold833/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 hold888/X hold888/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 hold877/X hold877/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13623__740 VPWR VGND VPWR VGND _14963_/CLK clkload34/A sky130_fd_sc_hd__inv_2
Xhold866 hold866/X hold866/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ VPWR VGND VGND VPWR _09986_/B _09984_/B _15608_/D sky130_fd_sc_hd__nor2_1
Xhold899 hold899/X hold899/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08935_ VPWR VGND _09869_/A _08935_/B _08935_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_29_203 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08866_ VPWR VGND VGND VPWR _08866_/X _15159_/Q _08918_/B sky130_fd_sc_hd__or2_1
X_07817_ VPWR VGND VGND VPWR _07817_/A _07900_/A _07878_/B sky130_fd_sc_hd__nor2_1
X_08797_ VGND VPWR VPWR VGND _15212_/D fanout35/X _08806_/S hold550/X sky130_fd_sc_hd__mux2_1
X_07748_ VGND VPWR _07748_/X _15598_/Q _15551_/Q _07751_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_38_792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07679_ VGND VPWR _07679_/B _07679_/Y _07679_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_10690_ VGND VPWR VGND VPWR _10690_/X _10697_/B1 _10685_/X _10689_/X _10469_/S sky130_fd_sc_hd__o211a_1
X_13472__589 VPWR VGND VPWR VGND _14747_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_09418_ _14634_/D fanout94/X fanout90/X _09416_/Y _09417_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09349_ VGND VPWR VPWR VGND _14697_/D hold709/X _09357_/S fanout86/X sky130_fd_sc_hd__mux2_1
X_12360_ VGND VPWR VGND VPWR _12360_/X _12863_/A1 _12355_/X _12359_/X _12472_/S sky130_fd_sc_hd__o211a_1
X_11311_ VPWR VGND VGND VPWR _11421_/C _14833_/Q _11408_/A sky130_fd_sc_hd__nand2_2
X_12291_ VGND VPWR VPWR VGND _12291_/X _12290_/X _12698_/S _12289_/X sky130_fd_sc_hd__mux2_1
X_11242_ VPWR VGND VGND VPWR _11242_/X _11250_/S _11242_/B sky130_fd_sc_hd__or2_1
XFILLER_5_858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13366__483 VPWR VGND VPWR VGND _14641_/CLK clkload51/A sky130_fd_sc_hd__inv_2
XFILLER_10_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11173_ VPWR VGND VGND VPWR _11173_/A _11173_/B _11173_/Y sky130_fd_sc_hd__nor2_1
X_10124_ VPWR VGND VGND VPWR _10124_/X _10615_/S _10124_/B sky130_fd_sc_hd__or2_1
XFILLER_76_832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14932_ _14932_/Q clkload29/A _14932_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10055_ VGND VPWR VGND VPWR _15639_/D _10060_/A _14801_/Q _12878_/B _08571_/B sky130_fd_sc_hd__o211a_1
XFILLER_48_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14863_ _14863_/Q _14863_/CLK _14863_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14794_ hold641/A _14794_/CLK _14794_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10957_ VGND VPWR VPWR VGND _10957_/X _14885_/Q _11179_/S hold425/A sky130_fd_sc_hd__mux2_1
X_10888_ VPWR VGND VGND VPWR _10888_/X _11110_/A _10888_/B sky130_fd_sc_hd__or2_1
X_12627_ VGND VPWR VPWR VGND _12627_/X _14890_/Q _12635_/B hold363/A sky130_fd_sc_hd__mux2_1
X_15415_ hold591/A _15415_/CLK _15415_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15346_ _15346_/Q _15346_/CLK _15346_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12558_ VGND VPWR VGND VPWR _12558_/X _15025_/Q _12743_/A2 _12735_/S _12557_/X sky130_fd_sc_hd__o211a_1
X_11509_ VGND VPWR VPWR VGND _11509_/X _11508_/X _11537_/S _15467_/Q sky130_fd_sc_hd__mux2_1
X_15277_ hold872/A _15277_/CLK _15277_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13607__724 VPWR VGND VPWR VGND _14947_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_12489_ VGND VPWR VGND VPWR _12489_/X _12486_/X _12488_/X _12489_/A1 _12722_/A1 sky130_fd_sc_hd__a211o_1
X_14228_ hold338/A _14228_/CLK _14228_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout609 VPWR VGND _08300_/S _08267_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_14159_ hold731/A _14159_/CLK _14159_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14189__907 _14189_/D _14189__907/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_39_512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08720_ VPWR VGND VPWR VGND _15272_/Q _08523_/B _08720_/X _08728_/B1 _14384_/Q _08722_/C1
+ sky130_fd_sc_hd__a221o_1
X_08651_ VPWR VGND VGND VPWR _08650_/X _08690_/S _08194_/Y _14406_/Q _08651_/X _08649_/X
+ sky130_fd_sc_hd__o221a_1
X_07602_ _15544_/D _07133_/Y fanout93/X fanout89/X _07601_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08582_ VPWR VGND VGND VPWR _08582_/A _08989_/B _08582_/Y sky130_fd_sc_hd__nor2_1
X_07533_ VPWR VGND VPWR VGND _07533_/X _07523_/B _07532_/Y _07531_/X _07527_/X _07523_/Y
+ sky130_fd_sc_hd__o32a_1
XFILLER_39_1424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07464_ VPWR VGND VGND VPWR _15450_/Q _08608_/B _15595_/Q sky130_fd_sc_hd__nand2_1
XFILLER_39_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14046__1163 VPWR VGND VPWR VGND _15418_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_09203_ VGND VPWR VPWR VGND _14890_/D hold1074/X _09213_/S clone146/X sky130_fd_sc_hd__mux2_1
X_07395_ VGND VPWR VGND VPWR _07395_/X _07855_/B _07859_/A _07819_/A sky130_fd_sc_hd__a21bo_1
X_09134_ VGND VPWR VPWR VGND _14964_/D fanout80/X _09157_/S hold813/X sky130_fd_sc_hd__mux2_1
X_13053__170 VPWR VGND VPWR VGND _14296_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_09065_ VGND VPWR VPWR VGND _15028_/D hold1047/X _09090_/S fanout80/X sky130_fd_sc_hd__mux2_1
Xhold630 hold630/X hold630/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08016_ VPWR VGND VPWR VGND clone20/X _15346_/Q clone13/X _08016_/X _15151_/Q sky130_fd_sc_hd__a22o_1
Xhold652 hold652/X hold652/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 hold663/X hold663/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 hold641/X hold641/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13975__1092 VPWR VGND VPWR VGND _15347_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
Xhold685 hold685/X hold685/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/X hold674/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 hold696/X hold696/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ VGND VPWR _07421_/Y _07563_/B _09967_/Y _10059_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_08918_ VPWR VGND VGND VPWR _08918_/X _15133_/Q _08918_/B sky130_fd_sc_hd__or2_1
XFILLER_40_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09898_ VPWR VGND VPWR VGND _09897_/X _08858_/Y _09893_/Y _14144_/D hold1145/X sky130_fd_sc_hd__a22o_1
Xhold1352 hold1352/X _14126_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13400__517 VPWR VGND VPWR VGND _14675_/CLK clkload20/A sky130_fd_sc_hd__inv_2
Xhold1330 _10051_/A _15637_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1341 _10044_/A _15634_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_1049 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1385 hold1385/X _14442_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 _09766_/A _14282_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1374 _09417_/A _14634_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08849_ VGND VPWR VPWR VGND _15164_/D _09692_/A0 _08850_/S hold498/X sky130_fd_sc_hd__mux2_1
Xhold1396 _08415_/B _14806_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11860_ VGND VPWR VGND VPWR _11860_/X _11859_/X _11858_/X _12119_/A1 _12017_/C1 sky130_fd_sc_hd__a211o_1
X_11791_ VGND VPWR VPWR VGND _11791_/X hold912/A _12589_/S hold551/A sky130_fd_sc_hd__mux2_1
X_10811_ VGND VPWR VPWR VGND _10811_/X _15018_/Q _11223_/S hold891/A sky130_fd_sc_hd__mux2_1
X_10742_ VGND VPWR VPWR VGND _10742_/X hold646/A _10742_/S hold595/A sky130_fd_sc_hd__mux2_1
X_15200_ hold404/A _15200_/CLK _15200_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10673_ VPWR VGND VPWR VGND _10672_/X _10729_/A _11973_/B _10673_/X sky130_fd_sc_hd__a21o_1
X_12412_ VGND VPWR VPWR VGND _12412_/X hold428/A _12726_/S hold688/A sky130_fd_sc_hd__mux2_1
X_12343_ VPWR VGND VPWR VGND _12342_/X _12473_/A _12602_/B1 _12343_/X sky130_fd_sc_hd__a21o_1
X_15131_ _15131_/Q _15131_/CLK _15131_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12274_ VGND VPWR VPWR VGND _12274_/X hold490/A _12689_/S hold207/A sky130_fd_sc_hd__mux2_1
X_15062_ _15062_/Q _15062_/CLK _15062_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11225_ VGND VPWR VGND VPWR _11225_/X _15029_/Q _11262_/A2 _11224_/X _10851_/A sky130_fd_sc_hd__o211a_1
XFILLER_67_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11156_ VGND VPWR VPWR VGND _11160_/B _14632_/Q _11179_/S _14664_/Q sky130_fd_sc_hd__mux2_1
X_11087_ VGND VPWR VPWR VGND _11087_/X _14566_/Q _11093_/S _14598_/Q sky130_fd_sc_hd__mux2_1
X_10107_ VGND VPWR VGND VPWR _10107_/X _10106_/X _10105_/X _10144_/S _10614_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_76_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14915_ _14915_/Q _14915_/CLK _14915_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10038_ VGND VPWR _10042_/B _15632_/Q _15631_/Q _10038_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_75_172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_64_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_64_846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14846_ _14846_/Q clkload20/A _14846_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14777_ hold357/A _14777_/CLK _14777_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11989_ VGND VPWR VPWR VGND _11989_/X _11986_/X _11995_/S _11985_/X sky130_fd_sc_hd__mux2_1
X_13999__1116 VPWR VGND VPWR VGND _15371_/CLK clkload11/A sky130_fd_sc_hd__inv_2
XFILLER_73_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07180_ _07972_/A _15462_/Q _07180_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_13037__154 VPWR VGND VPWR VGND _14280_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_15329_ _15329_/Q _15329_/CLK _15329_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12965__82 VPWR VGND VPWR VGND _14208_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_13841__958 VPWR VGND VPWR VGND _15213_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
Xfanout439 VGND VPWR _11096_/C1 _11218_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout417 VGND VPWR fanout424/X _12868_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout428 VGND VPWR _10706_/C1 _10693_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09821_ VGND VPWR VPWR VGND _14231_/D fanout16/X _09833_/S hold175/X sky130_fd_sc_hd__mux2_1
X_13694__811 VPWR VGND VPWR VGND _15034_/CLK clkload37/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09752_ VGND VPWR VPWR VGND _14294_/D fanout12/X _09763_/S hold410/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08703_ VGND VPWR VGND VPWR _08703_/X _08714_/A2 _08722_/C1 hold1438/X _08702_/X
+ sky130_fd_sc_hd__a211o_1
X_13735__852 VPWR VGND VPWR VGND _15107_/CLK clkload30/A sky130_fd_sc_hd__inv_2
XFILLER_67_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09683_ VGND VPWR VPWR VGND _14357_/D hold929/X _09693_/S fanout9/A sky130_fd_sc_hd__mux2_1
X_08634_ VGND VPWR VGND VPWR _08700_/A2 _14385_/Q _08194_/B _08634_/X sky130_fd_sc_hd__o21ba_1
X_08565_ VPWR VGND VGND VPWR _15555_/Q _08565_/Y _08591_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07516_ VGND VPWR VGND VPWR _07539_/B _07547_/B _07547_/C _07547_/A _07515_/Y sky130_fd_sc_hd__a211o_1
Xfanout13 VGND VPWR _08091_/X fanout13/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_08496_ VPWR VGND VPWR VGND _08500_/B _09912_/A _09937_/B _08507_/C sky130_fd_sc_hd__a21oi_1
Xfanout46 VGND VPWR _07910_/X fanout46/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout35 VGND VPWR fanout36/X fanout35/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout24 VPWR VGND fanout24/X _08032_/X VPWR VGND sky130_fd_sc_hd__buf_6
X_07447_ VPWR VGND VGND VPWR _07447_/A _08575_/A _07447_/B sky130_fd_sc_hd__nand2_1
Xfanout68 VPWR VGND fanout68/X fanout71/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout57 VPWR VGND VGND VPWR clone55/A fanout57/X sky130_fd_sc_hd__buf_8
Xfanout79 VPWR VGND VGND VPWR _07643_/X fanout79/X sky130_fd_sc_hd__buf_8
XFILLER_22_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07378_ VPWR VGND _08064_/B _08081_/B _08081_/A _07356_/Y _07357_/Y VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_10_459 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09117_ VGND VPWR VPWR VGND _14978_/D hold343/X _09128_/S fanout13/X sky130_fd_sc_hd__mux2_1
X_09048_ VGND VPWR VPWR VGND _15042_/D hold796/X _09059_/S fanout14/X sky130_fd_sc_hd__mux2_1
Xhold471 hold471/X hold471/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 hold460/X hold460/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_916 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold493 hold493/X hold493/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 hold482/X hold482/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ VGND VPWR VPWR VGND _11010_/X hold662/A _11165_/S hold289/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1160 hold1160/X _11553_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1193 hold1193/X _15333_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 hold1171/X _15154_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13478__595 VPWR VGND VPWR VGND _14753_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_2_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14700_ hold648/A _14700_/CLK _14700_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11912_ VGND VPWR VPWR VGND _11912_/X hold538/A _12205_/S hold312/A sky130_fd_sc_hd__mux2_1
Xhold1182 hold1182/X _14457_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11843_ VGND VPWR VPWR VGND _11844_/B _11842_/Y _12176_/S _11834_/Y sky130_fd_sc_hd__mux2_1
X_14631_ hold629/A _14631_/CLK _14631_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1207 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14562_ hold603/A _14562_/CLK _14562_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11774_ VPWR VGND VGND VPWR _11774_/X hold362/A _12006_/B sky130_fd_sc_hd__or2_1
X_14493_ _14493_/Q _14493_/CLK _14493_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10725_ VGND VPWR VGND VPWR _10725_/X _10745_/A1 _10721_/X _10724_/X _10741_/C1 sky130_fd_sc_hd__o211a_1
X_10656_ VPWR VGND VGND VPWR _10656_/X hold375/A _10664_/S sky130_fd_sc_hd__or2_1
Xclkload16 VGND VPWR VGND VPWR clkload16/Y clkload16/A sky130_fd_sc_hd__inv_8
X_15114_ hold543/A _15114_/CLK _15114_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkload49 clkload49/Y clkload49/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload27 clkload27/Y clkload27/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
Xclkload38 clkload38/Y clkload38/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
X_10587_ VGND VPWR VPWR VGND _10587_/X hold857/A _10730_/S hold634/A sky130_fd_sc_hd__mux2_1
X_12326_ VGND VPWR VPWR VGND _12326_/X hold785/A _12594_/B hold565/A sky130_fd_sc_hd__mux2_1
X_12257_ VPWR VGND VPWR VGND _12256_/X _12703_/A1 _12255_/X _12257_/X sky130_fd_sc_hd__a21o_1
X_15045_ hold736/A _15045_/CLK _15045_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11208_ VPWR VGND VPWR VGND _11207_/X _11218_/A1 _11206_/X _11208_/Y sky130_fd_sc_hd__a21oi_1
X_12188_ VGND VPWR VGND VPWR _12188_/X hold909/A _12188_/A2 _12180_/S _12187_/X sky130_fd_sc_hd__o211a_1
XFILLER_29_1445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14045__1162 VPWR VGND VPWR VGND _15417_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_11139_ VGND VPWR VPWR VGND _11139_/X _14963_/Q _11146_/B hold540/A sky130_fd_sc_hd__mux2_1
X_13719__836 VPWR VGND VPWR VGND _15059_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XFILLER_49_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_49_662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_37_802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_64_654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_64_621 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_868 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14829_ _14829_/Q clkload30/A _14829_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08350_ VGND VPWR VPWR VGND _15423_/D hold371/X _08356_/S fanout64/X sky130_fd_sc_hd__mux2_1
XFILLER_24_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13974__1091 VPWR VGND VPWR VGND _15346_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_07301_ VGND VPWR VGND VPWR _07311_/A _14400_/Q _07301_/A2 _07301_/B1 _15466_/Q sky130_fd_sc_hd__o211a_1
X_08281_ _08281_/X _08278_/X _08279_/X _08280_/X _08294_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07232_ VPWR VGND _08257_/B _08290_/B _08278_/A _15445_/Q _07226_/Y VGND VPWR sky130_fd_sc_hd__a31o_1
X_13271__388 VPWR VGND VPWR VGND _14546_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_07163_ VPWR VGND VPWR VGND _07639_/A _07163_/A _07640_/A sky130_fd_sc_hd__or2_2
X_07094_ VPWR VGND VPWR VGND _07369_/A _15450_/Q sky130_fd_sc_hd__inv_2
Xfanout214 VPWR VGND _12588_/A1 fanout217/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout203 VGND VPWR _12226_/A1 _12156_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout247 VGND VPWR _12666_/A1 _12740_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09804_ VGND VPWR VPWR VGND _14248_/D clone49/A _09827_/S hold276/X sky130_fd_sc_hd__mux2_1
Xfanout225 VGND VPWR _12863_/A1 _12485_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout236 VPWR VGND _12008_/C1 _12193_/C1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout258 _12139_/S _12213_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout269 VPWR VGND _12584_/A _07912_/X VPWR VGND sky130_fd_sc_hd__buf_4
X_07996_ VGND VPWR VPWR VGND _08198_/S _07597_/X _07996_/X _10058_/A1 sky130_fd_sc_hd__o21a_4
X_13165__282 VPWR VGND VPWR VGND _14440_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_09735_ VGND VPWR VPWR VGND _14311_/D _09757_/S fanout76/X hold1252/X sky130_fd_sc_hd__mux2_4
X_09666_ VGND VPWR VPWR VGND _14374_/D _09675_/S hold1240/X fanout72/X sky130_fd_sc_hd__mux2_4
XFILLER_76_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08617_ VPWR VGND VGND VPWR _08617_/A _09010_/B _08617_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_676 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09597_ VGND VPWR VPWR VGND _14471_/D fanout78/X _09619_/S hold582/X sky130_fd_sc_hd__mux2_1
X_08548_ VPWR VGND VPWR VGND _08548_/B _08548_/C _08548_/A _08548_/X sky130_fd_sc_hd__or3_1
X_13512__629 VPWR VGND VPWR VGND _14787_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_08479_ VGND VPWR VGND VPWR _08479_/X hold1217/X _08483_/A2 _08478_/X _11431_/C1
+ sky130_fd_sc_hd__o211a_1
X_11490_ VGND VPWR VPWR VGND _11490_/X _15082_/Q _11490_/S _15080_/Q sky130_fd_sc_hd__mux2_1
X_10510_ VGND VPWR VPWR VGND _10510_/X _10509_/X _10510_/S _10508_/X sky130_fd_sc_hd__mux2_1
X_10441_ VGND VPWR VPWR VGND _10441_/X _15008_/Q _10554_/S hold678/A sky130_fd_sc_hd__mux2_1
X_13863__980 VPWR VGND VPWR VGND _15235_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_10372_ VGND VPWR VPWR VGND _10372_/X hold562/A _10702_/S hold747/A sky130_fd_sc_hd__mux2_1
XFILLER_3_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12111_ VGND VPWR VGND VPWR _12111_/X _12193_/C1 _12106_/X _12110_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
X_12042_ VGND VPWR VPWR VGND _12042_/X hold417/A _12043_/B hold402/A sky130_fd_sc_hd__mux2_1
X_13406__523 VPWR VGND VPWR VGND _14681_/CLK clkload7/A sky130_fd_sc_hd__inv_2
Xhold290 hold290/X hold290/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13998__1115 VPWR VGND VPWR VGND _15370_/CLK clkload35/A sky130_fd_sc_hd__inv_2
Xfanout792 VGND VPWR fanout802/X _09912_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout770 VGND VPWR _08104_/B _07972_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout781 VPWR VGND _07265_/B1 _07144_/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12875_ VGND VPWR VPWR VGND _15599_/D _07616_/X _14802_/D _15599_/Q sky130_fd_sc_hd__mux2_1
XFILLER_57_1162 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11826_ VPWR VGND VGND VPWR _11807_/Y _11825_/X _12269_/B _15451_/Q _15451_/D _11341_/A
+ sky130_fd_sc_hd__o221a_1
X_15594_ _15594_/Q clkload50/A _15594_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14614_ hold916/A _14614_/CLK _14614_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14545_ _14545_/Q _14545_/CLK _14545_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11757_ VPWR VGND VGND VPWR _11757_/X _12098_/A _11757_/B sky130_fd_sc_hd__or2_1
X_10708_ VPWR VGND _10708_/X _10698_/X _10694_/X _10737_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
X_11688_ VGND VPWR VPWR VGND _11688_/X hold492/A _12052_/S hold259/A sky130_fd_sc_hd__mux2_1
X_14476_ _14476_/Q _14476_/CLK _14476_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10639_ VGND VPWR VPWR VGND _10639_/X hold996/A _10720_/S hold533/A sky130_fd_sc_hd__mux2_1
X_12309_ VGND VPWR VPWR VGND _12309_/X hold847/A _12577_/S hold767/A sky130_fd_sc_hd__mux2_1
X_12935__52 VPWR VGND VPWR VGND _14178_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_13149__266 VPWR VGND VPWR VGND _14424_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_15028_ _15028_/Q _15028_/CLK _15028_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_69_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07850_ VGND VPWR VPWR VGND _15536_/D clone55/A _08231_/S hold162/X sky130_fd_sc_hd__mux2_1
X_07781_ VPWR VGND VPWR VGND _08146_/B _07750_/B _07748_/X _08126_/A sky130_fd_sc_hd__a21o_1
XFILLER_42_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 VGND VPWR input3/X ui_in[1] VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_09520_ VGND VPWR VPWR VGND _14539_/D fanout95/X _09520_/S hold803/X sky130_fd_sc_hd__mux2_1
X_09451_ VPWR VGND _09834_/A _09451_/X _09486_/C VPWR VGND sky130_fd_sc_hd__and2_2
XFILLER_80_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_40_819 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08402_ VGND VPWR VPWR VGND _15375_/D fanout5/X _08411_/S hold765/X sky130_fd_sc_hd__mux2_1
X_09382_ VPWR VGND VGND VPWR hold1365/X _09411_/S _09382_/Y sky130_fd_sc_hd__nand2b_1
X_08333_ VGND VPWR VPWR VGND _15486_/D _09550_/A1 _08338_/S hold958/X sky130_fd_sc_hd__mux2_1
X_08264_ VGND VPWR _08263_/X _08294_/B1 _08264_/Y _08260_/X VPWR VGND sky130_fd_sc_hd__o21ai_1
X_13847__964 VPWR VGND VPWR VGND _15219_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_08195_ VPWR VGND VPWR VGND _08232_/B _08195_/C _08195_/A _08195_/X sky130_fd_sc_hd__or3_1
X_07215_ VGND VPWR VPWR VGND _07220_/S _15594_/Q _14383_/Q _12845_/A sky130_fd_sc_hd__mux2_2
X_07146_ VGND VPWR _07304_/A2 _07304_/B1 _07149_/B _14410_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_10_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_74_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07979_ VPWR VGND VPWR VGND _15137_/Q clone19/X _15348_/Q _07558_/B _07979_/X sky130_fd_sc_hd__a22o_2
X_09718_ VGND VPWR VPWR VGND _14325_/D fanout9/X _09728_/S hold717/X sky130_fd_sc_hd__mux2_1
X_10990_ VGND VPWR VGND VPWR _10990_/X hold964/A _11003_/A2 _10989_/X _10995_/S sky130_fd_sc_hd__o211a_1
X_09649_ VGND VPWR VPWR VGND _14421_/D hold766/X _09659_/S fanout10/X sky130_fd_sc_hd__mux2_1
XFILLER_55_484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_35_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12660_ VGND VPWR VGND VPWR _12660_/X _14891_/Q _12669_/A2 _12655_/S _12659_/X sky130_fd_sc_hd__o211a_1
X_11611_ VGND VPWR VPWR VGND _11611_/X _11608_/X _12100_/S _11607_/X sky130_fd_sc_hd__mux2_1
X_12591_ VGND VPWR VPWR VGND _12591_/X _12590_/X _12591_/S _12589_/X sky130_fd_sc_hd__mux2_1
X_14044__1161 VPWR VGND VPWR VGND _15416_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_14330_ hold700/A _14330_/CLK _14330_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11542_ VGND VPWR VPWR VGND _11542_/B _11269_/B _11542_/A _15431_/D sky130_fd_sc_hd__or3b_1
XFILLER_11_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14261_ hold901/A _14261_/CLK _14261_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11473_ VGND VPWR VPWR VGND _11473_/X _11472_/X _11476_/S _15455_/Q sky130_fd_sc_hd__mux2_1
X_14192_ _14192_/Q _14192_/CLK _14192_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10424_ VGND VPWR VPWR VGND _10424_/X _14196_/Q _10743_/B hold303/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10355_ VGND VPWR VGND VPWR _10355_/X _10698_/A1 _10351_/X _10354_/X _10697_/B1 sky130_fd_sc_hd__o211a_1
XFILLER_65_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13640__757 VPWR VGND VPWR VGND _14980_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_10286_ VGND VPWR VPWR VGND _10286_/X hold816/A _10670_/S hold671/A sky130_fd_sc_hd__mux2_1
X_13973__1090 VPWR VGND VPWR VGND _15345_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_12025_ VGND VPWR VGND VPWR _12025_/X _11894_/S _12021_/X _12024_/X _12189_/C1 sky130_fd_sc_hd__o211a_1
X_13493__610 VPWR VGND VPWR VGND _14768_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_73_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12858_ VGND VPWR VPWR VGND _15582_/D _08053_/X _12860_/S _08286_/B sky130_fd_sc_hd__mux2_1
X_13534__651 VPWR VGND VPWR VGND _14865_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_11809_ VGND VPWR VPWR VGND _11809_/X hold859/A _12747_/S hold491/A sky130_fd_sc_hd__mux2_1
X_15577_ _15577_/Q clkload32/A _15577_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12789_ VPWR VGND VGND VPWR _12789_/A _12789_/Y _12789_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_381 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14528_ _14528_/Q _14528_/CLK _14528_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14459_ hold694/A _14459_/CLK _14459_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_72_Right_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08951_ VPWR VGND VGND VPWR _08936_/X hold1011/X _08933_/Y _15120_/Q _08951_/X _11567_/A
+ sky130_fd_sc_hd__o221a_1
X_08882_ VPWR VGND VGND VPWR _08882_/X _08882_/A _08926_/B sky130_fd_sc_hd__or2_1
X_07902_ VGND VPWR VPWR VGND _07902_/X _15085_/Q _10072_/B _07307_/B _07972_/B sky130_fd_sc_hd__o2bb2a_1
X_07833_ VPWR VGND _08145_/A _08155_/A _15551_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_42_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07764_ VGND VPWR VPWR VGND _15574_/Q _12855_/A0 _07765_/B _07769_/B sky130_fd_sc_hd__or3b_1
XFILLER_38_952 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_77_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07695_ VGND VPWR VPWR VGND _07695_/X _10066_/A _07857_/A _07693_/Y sky130_fd_sc_hd__mux2_1
X_09503_ VGND VPWR VPWR VGND _14556_/D fanout35/X _09513_/S hold584/X sky130_fd_sc_hd__mux2_1
XFILLER_77_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09434_ VGND VPWR VPWR VGND _14618_/D fanout28/X _09441_/S hold515/X sky130_fd_sc_hd__mux2_1
X_13277__394 VPWR VGND VPWR VGND _14552_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_09365_ VGND VPWR VPWR VGND _14681_/D hold440/X _09379_/S fanout25/X sky130_fd_sc_hd__mux2_1
XFILLER_21_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_30 _14408_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08316_ VGND VPWR VPWR VGND _15503_/D clone5/A _08318_/S hold1077/X sky130_fd_sc_hd__mux2_1
X_13997__1114 VPWR VGND VPWR VGND _15369_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XANTENNA_41 _12866_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_09296_ VGND VPWR VPWR VGND _14745_/D _09310_/S fanout23/X hold1201/X sky130_fd_sc_hd__mux2_4
X_08247_ VGND VPWR VPWR VGND _08247_/A _08247_/X _08247_/B sky130_fd_sc_hd__xor2_1
XANTENNA_63 _09272_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_74 _09756_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_384 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_52 _10505_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_96 fanout234/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_85 _08780_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08178_ VPWR VGND VGND VPWR _08178_/A1 _08172_/X _08177_/X _08178_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_1426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_723 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10140_ VGND VPWR VPWR VGND _10140_/X hold873/A _10140_/S hold483/A sky130_fd_sc_hd__mux2_1
X_10071_ VGND VPWR _10071_/X _10071_/B _10071_/A _10071_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_43_1058 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13518__635 VPWR VGND VPWR VGND _14793_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_6_Left_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10973_ VGND VPWR VPWR VGND _10973_/X hold482/A _10994_/S hold313/A sky130_fd_sc_hd__mux2_1
X_15500_ hold881/A _15500_/CLK _15500_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_955 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12712_ VPWR VGND _12712_/X _12711_/X _12707_/X _12694_/S _12703_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15431_ _15431_/Q clkload47/A _15431_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12643_ VGND VPWR VPWR VGND _12643_/X _14344_/Q _12651_/S hold247/A sky130_fd_sc_hd__mux2_1
X_12574_ VPWR VGND VPWR VGND _12573_/X _12703_/A1 _12572_/X _12574_/Y sky130_fd_sc_hd__a21oi_1
X_15362_ _15362_/Q _15362_/CLK _15362_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14313_ hold323/A _14313_/CLK _14313_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15293_ hold883/A _15293_/CLK _15293_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11525_ VGND VPWR VPWR VGND _15092_/D _11524_/X _11528_/S hold1422/X sky130_fd_sc_hd__mux2_1
XFILLER_7_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14244_ hold364/A _14244_/CLK _14244_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13070__187 VPWR VGND VPWR VGND _14313_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_11456_ VGND VPWR VPWR VGND _15069_/D _11455_/X _11480_/S hold1361/X sky130_fd_sc_hd__mux2_1
X_12905__22 VPWR VGND VPWR VGND _14147_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_14175_ hold767/A _14175_/CLK _14175_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11387_ VGND VPWR VPWR VGND _11387_/X _11386_/X _11387_/S _14850_/Q sky130_fd_sc_hd__mux2_1
X_10407_ VGND VPWR VGND VPWR _10407_/X hold821/A _10688_/A2 _10406_/X _10703_/A sky130_fd_sc_hd__o211a_1
X_10338_ VPWR VGND _10338_/X _10328_/X _10324_/X _11218_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_79_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10269_ VGND VPWR VPWR VGND _10269_/X hold864/A _10609_/S hold395/A sky130_fd_sc_hd__mux2_1
X_12008_ VGND VPWR VGND VPWR _12008_/X _12005_/X _12007_/X _12008_/A1 _12008_/C1 sky130_fd_sc_hd__a211o_1
X_07480_ VPWR VGND VGND VPWR _07573_/A _07564_/B _07480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15629_ _15629_/Q clkload49/A _15629_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09150_ VGND VPWR VPWR VGND _14948_/D fanout21/X _09161_/S hold894/X sky130_fd_sc_hd__mux2_1
X_08101_ VPWR VGND VGND VPWR _08277_/S _08101_/Y _12783_/B sky130_fd_sc_hd__nand2_1
X_09081_ VGND VPWR VPWR VGND _15012_/D hold1078/X _09091_/S fanout21/X sky130_fd_sc_hd__mux2_1
X_13311__428 VPWR VGND VPWR VGND _14586_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_08032_ VGND VPWR VGND VPWR _08032_/X _08024_/X _08032_/C _08032_/B _08032_/A sky130_fd_sc_hd__or4b_4
Xhold812 hold812/X hold812/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold801 hold801/X hold801/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 hold823/X hold823/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 hold845/X hold845/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 hold834/X hold834/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/X hold867/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ VPWR VGND VPWR VGND _15607_/Q hold807/A hold1314/X _09983_/Y sky130_fd_sc_hd__a21oi_1
Xhold889 hold889/X hold889/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold878 hold878/X hold878/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 hold856/X hold856/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ VPWR VGND VPWR VGND _09970_/B _15162_/Q _09906_/A _08935_/B sky130_fd_sc_hd__a21o_1
X_08865_ VGND VPWR VGND VPWR _08865_/X hold1257/X _08893_/A2 _08864_/X _09024_/A sky130_fd_sc_hd__o211a_1
X_13205__322 VPWR VGND VPWR VGND _14480_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_14043__1160 VPWR VGND VPWR VGND _15415_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_08796_ VGND VPWR VPWR VGND _15213_/D fanout40/X _08811_/S hold277/X sky130_fd_sc_hd__mux2_1
X_07816_ VGND VPWR VGND VPWR _07900_/A _07387_/X _07351_/Y _07899_/A sky130_fd_sc_hd__a21bo_1
XFILLER_77_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07747_ VGND VPWR _07747_/X _15599_/Q _15552_/Q _07751_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_41_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07678_ VPWR VGND VPWR VGND _07694_/A _07693_/A _07316_/A _07679_/B sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09417_ VPWR VGND VGND VPWR _09417_/X _09417_/A _09446_/S sky130_fd_sc_hd__or2_1
X_09348_ _14698_/D fanout91/X fanout87/X _09357_/S _09347_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_32_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11310_ VPWR VGND VPWR VGND _14831_/Q _14829_/Q _14830_/Q _14832_/Q _11421_/B sky130_fd_sc_hd__or4_2
X_09279_ _14762_/D fanout92/X fanout88/X _09277_/Y _09278_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_12290_ VGND VPWR VPWR VGND _12290_/X hold852/A _12701_/S hold762/A sky130_fd_sc_hd__mux2_1
X_11241_ VGND VPWR VPWR VGND _11241_/X _14474_/Q _11241_/S _14762_/Q sky130_fd_sc_hd__mux2_1
XFILLER_10_1057 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11172_ VGND VPWR VPWR VGND _11173_/B _11171_/Y _11246_/S _11163_/Y sky130_fd_sc_hd__mux2_1
XFILLER_79_137 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10123_ VGND VPWR VPWR VGND _10123_/X hold647/A _10353_/S hold342/A sky130_fd_sc_hd__mux2_1
X_14931_ _14931_/Q clkload29/A _14931_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10054_ VPWR VGND VGND VPWR _11340_/A _11973_/B _10054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14862_ hold860/A _14862_/CLK _14862_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13752__869 VPWR VGND VPWR VGND _15124_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_14793_ hold560/A _14793_/CLK _14793_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10956_ VGND VPWR VGND VPWR _10956_/X hold961/A _11184_/A2 _10955_/X _11178_/C1 sky130_fd_sc_hd__o211a_1
X_10887_ VGND VPWR VPWR VGND _10890_/B _15502_/Q _11109_/S _14528_/Q sky130_fd_sc_hd__mux2_1
XFILLER_32_958 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15414_ hold380/A _15414_/CLK _15414_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_969 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12626_ VGND VPWR VGND VPWR _12626_/X _14963_/Q _12743_/A2 _12737_/B1 _12625_/X sky130_fd_sc_hd__o211a_1
X_15345_ _15345_/Q _15345_/CLK _15345_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12557_ VPWR VGND VGND VPWR _12557_/X hold332/A _12671_/S sky130_fd_sc_hd__or2_1
X_13646__763 VPWR VGND VPWR VGND _14986_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_11508_ VGND VPWR VPWR VGND _11508_/X _15088_/Q _11535_/C _15086_/Q sky130_fd_sc_hd__mux2_1
X_15276_ hold982/A _15276_/CLK _15276_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_8_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12488_ VGND VPWR VGND VPWR _12488_/X _15023_/Q _12488_/A2 _12470_/S _12487_/X sky130_fd_sc_hd__o211a_1
X_11439_ VGND VPWR VGND VPWR _14934_/D _14822_/Q _11439_/A2 _11438_/X _11347_/A sky130_fd_sc_hd__o211a_1
X_14227_ hold197/A _14227_/CLK _14227_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14158_ hold439/A _14158_/CLK _14158_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1378 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13996__1113 VPWR VGND VPWR VGND _15368_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_08650_ VPWR VGND VGND VPWR _08650_/X _14390_/Q _08664_/B sky130_fd_sc_hd__or2_1
X_07601_ VPWR VGND VGND VPWR _07601_/X _07601_/A _08231_/S sky130_fd_sc_hd__or2_1
XFILLER_78_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08581_ VGND VPWR VPWR VGND _08989_/B _15553_/Q _08591_/B _10060_/C _08580_/Y sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_281 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07532_ VPWR VGND VPWR VGND _07531_/A _07531_/C _07531_/B _07532_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_1436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07463_ VPWR VGND VGND VPWR _15450_/Q _15595_/Q _07489_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09202_ VGND VPWR VPWR VGND _09213_/S hold1226/X clone49/X _14891_/D sky130_fd_sc_hd__mux2_2
X_13952__1069 VPWR VGND VPWR VGND _15324_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_09133_ VGND VPWR VPWR VGND _14965_/D fanout83/X _09157_/S hold932/X sky130_fd_sc_hd__mux2_1
X_07394_ VPWR VGND VPWR VGND _07300_/B _15466_/Q _07878_/A _07855_/B sky130_fd_sc_hd__a21o_1
X_09064_ VGND VPWR VPWR VGND _15029_/D hold1103/X _09088_/S fanout83/X sky130_fd_sc_hd__mux2_1
Xhold620 hold620/X hold620/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08015_ VGND VPWR VPWR VGND _15528_/D _08014_/X _08300_/S hold166/X sky130_fd_sc_hd__mux2_1
Xhold653 hold653/X hold653/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 hold642/X hold642/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 hold631/X hold631/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 hold697/X hold697/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 hold686/X hold686/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold664 hold664/X hold664/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 hold675/X hold675/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12896__13 VPWR VGND VPWR VGND _14138_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_09966_ VGND VPWR VPWR VGND _15260_/Q _10053_/B _11458_/S _09966_/X sky130_fd_sc_hd__or3b_1
X_14213__931 _14213_/D _14213__931/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09897_ VPWR VGND VPWR VGND _08859_/C _15480_/Q _09907_/S _09897_/X sky130_fd_sc_hd__a21o_1
X_08917_ VGND VPWR VGND VPWR _15134_/D hold1328/X _08919_/A2 _08916_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
X_08848_ VGND VPWR VPWR VGND _15165_/D _09229_/A0 _08850_/S hold984/X sky130_fd_sc_hd__mux2_1
Xhold1342 hold1342/X _15614_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1331 _15637_/D _10051_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1320 hold1320/X _15611_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 hold1364/X _15142_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 hold1386/X _15070_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 hold1375/X _15291_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1353 _09453_/A _14602_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1397 _08306_/A _15512_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08779_ VGND VPWR VPWR VGND _15227_/D fanout95/X _08779_/S hold160/X sky130_fd_sc_hd__mux2_1
X_11790_ VGND VPWR VPWR VGND _11794_/B hold374/A _12589_/S hold606/A sky130_fd_sc_hd__mux2_1
X_10810_ VGND VPWR VPWR VGND _10814_/B hold853/A _11223_/S hold663/A sky130_fd_sc_hd__mux2_1
X_13589__706 VPWR VGND VPWR VGND _14920_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_10741_ VGND VPWR VGND VPWR _10741_/X _10738_/X _10740_/X _10745_/A1 _10741_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_41_755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_55_1293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13333__450 VPWR VGND VPWR VGND _14608_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_10672_ VPWR VGND _10672_/X _10671_/X _10667_/X _10728_/S _10663_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_16_1222 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12411_ VGND VPWR VGND VPWR _12411_/X _12408_/X _12410_/X _12737_/B1 _12739_/C1 sky130_fd_sc_hd__a211o_1
Xclone20 VGND VPWR clone20/X clone20/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_20_clk _14821_/CLK clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_12_1119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12342_ VPWR VGND _12342_/X _12341_/X _12337_/X _12583_/S _12333_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15130_ _15130_/Q _15130_/CLK _15130_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12273_ VGND VPWR VPWR VGND _12273_/X _14334_/Q _12282_/S hold321/A sky130_fd_sc_hd__mux2_1
X_15061_ hold509/A _15061_/CLK _15061_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11224_ VPWR VGND VGND VPWR _11224_/X hold359/A _11261_/B sky130_fd_sc_hd__or2_1
XFILLER_4_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11155_ VPWR VGND VGND VPWR _11136_/Y _11154_/X _12677_/A2 _14407_/Q _14407_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_11086_ VGND VPWR VGND VPWR _11086_/X _14342_/Q _11262_/A2 _11085_/X _11086_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_0_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10106_ VGND VPWR VPWR VGND _10106_/X hold860/A _10609_/S hold517/A sky130_fd_sc_hd__mux2_1
X_14914_ hold387/A _14914_/CLK _14914_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10037_ VGND VPWR VPWR VGND _10037_/A _15631_/D _10038_/C sky130_fd_sc_hd__xor2_1
X_13182__299 VPWR VGND VPWR VGND _14457_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_48_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14845_ _14845_/Q clkload20/A _14845_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14776_ hold811/A _14776_/CLK _14776_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11988_ VGND VPWR VGND VPWR _11988_/X _12008_/A1 _11984_/X _11987_/X _12017_/C1 sky130_fd_sc_hd__o211a_1
X_10939_ VGND VPWR VGND VPWR _10939_/X _11178_/C1 _10935_/X _10938_/X _11180_/C1 sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_9_Left_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13076__193 VPWR VGND VPWR VGND _14319_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_73_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_clk clkload20/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12609_ VGND VPWR VGND VPWR _12609_/X _12737_/B1 _12605_/X _12608_/X _12739_/C1 sky130_fd_sc_hd__o211a_1
X_15328_ _15328_/Q _15328_/CLK _15328_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1399 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15259_ _15259_/Q _15259_/CLK _15259_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13880__997 VPWR VGND VPWR VGND _15252_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
Xfanout429 VGND VPWR _10505_/A1 _10706_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout418 VGND VPWR _11185_/C1 _11180_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09820_ VGND VPWR VPWR VGND _14232_/D fanout19/X _09825_/S hold302/X sky130_fd_sc_hd__mux2_1
X_12980__97 VPWR VGND VPWR VGND _14223_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
Xfanout407 VGND VPWR _10622_/C1 _10614_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09751_ VGND VPWR VPWR VGND _14295_/D fanout15/X _09763_/S hold227/X sky130_fd_sc_hd__mux2_1
X_08702_ VGND VPWR VGND VPWR _08702_/X _14391_/Q _08664_/B _08711_/B1 _08644_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13774__891 VPWR VGND VPWR VGND _15146_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_09682_ VGND VPWR VPWR VGND _14358_/D hold875/X _09693_/S fanout13/X sky130_fd_sc_hd__mux2_1
X_08633_ VGND VPWR VGND VPWR _15299_/D hold1354/X _08701_/A2 _08632_/X _12233_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08564_ VGND VPWR VGND VPWR _15313_/D hold905/X _08628_/A2 _08563_/X _11337_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_70_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07515_ VPWR VGND VPWR VGND _07515_/Y _07515_/A sky130_fd_sc_hd__inv_2
X_08495_ VPWR VGND VPWR VGND _08495_/A2 _15638_/Q _08493_/Y _08738_/B sky130_fd_sc_hd__a21o_1
X_13317__434 VPWR VGND VPWR VGND _14592_/CLK clkload45/A sky130_fd_sc_hd__inv_2
Xfanout47 VGND VPWR fanout47/X _07910_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout36 VGND VPWR _07976_/X fanout36/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout14 VPWR VGND fanout14/X _08091_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout25 VGND VPWR _08032_/X fanout25/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07446_ VPWR VGND VGND VPWR _15456_/Q _07447_/B _07714_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_1411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout69 VGND VPWR fanout71/X fanout69/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout58 VGND VPWR clone55/A fanout58/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07377_ VPWR VGND VPWR VGND _08117_/B _08117_/A _07376_/Y _08081_/B sky130_fd_sc_hd__a21oi_1
X_12990__107 VPWR VGND VPWR VGND _14233_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_09116_ VGND VPWR VPWR VGND _14979_/D hold899/X _09128_/S _08070_/X sky130_fd_sc_hd__mux2_1
X_09047_ VGND VPWR VPWR VGND _15043_/D hold402/X _09059_/S fanout17/X sky130_fd_sc_hd__mux2_1
Xhold472 hold472/X hold472/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold461/X hold461/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 hold450/X hold450/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 hold494/X hold494/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 hold483/X hold483/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09949_ VPWR VGND VGND VPWR _09954_/C _09949_/Y _09949_/B sky130_fd_sc_hd__nand2_1
Xhold1150 hold1150/X _15217_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1057 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1172 hold1172/X _14148_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 hold1183/X _14560_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 hold1161/X _15150_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_527 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11911_ VGND VPWR VPWR VGND _11911_/X _14196_/Q _12228_/B hold303/A sky130_fd_sc_hd__mux2_1
Xhold1194 hold1194/X _14376_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14630_ _14630_/Q _14630_/CLK _14630_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11842_ VPWR VGND VPWR VGND _11841_/X _12175_/A1 _11840_/X _11842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14561_ _14561_/Q _14561_/CLK _14561_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11773_ VGND VPWR VPWR VGND _11773_/X _11772_/X _12106_/S _11771_/X sky130_fd_sc_hd__mux2_1
X_10724_ VPWR VGND VGND VPWR _10724_/X _10732_/S _10724_/B sky130_fd_sc_hd__or2_1
X_14492_ hold974/A _14492_/CLK _14492_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10655_ VPWR VGND VGND VPWR _10729_/A _10655_/B _10655_/Y sky130_fd_sc_hd__nor2_1
X_13995__1112 VPWR VGND VPWR VGND _15367_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_6_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14022__1139 VPWR VGND VPWR VGND _15394_/CLK clkload34/A sky130_fd_sc_hd__inv_2
Xclkload17 VGND VPWR VPWR VGND clkload17/A clkload17/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload28 VPWR VGND VGND VPWR clkload28/Y clkload28/A sky130_fd_sc_hd__inv_16
X_15113_ hold791/A _15113_/CLK _15113_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12325_ VPWR VGND VGND VPWR _12584_/A _12325_/B _12325_/Y sky130_fd_sc_hd__nor2_1
Xclkload39 VGND VPWR VPWR VGND clkload39/A clkload39/Y sky130_fd_sc_hd__clkinv_4
X_10586_ VGND VPWR VPWR VGND _10586_/X hold898/A _10730_/S hold799/A sky130_fd_sc_hd__mux2_1
X_13110__227 VPWR VGND VPWR VGND _14353_/CLK clkload49/A sky130_fd_sc_hd__inv_2
X_12256_ VGND VPWR VPWR VGND _12256_/X _12251_/X _12256_/S _12250_/X sky130_fd_sc_hd__mux2_1
X_15044_ hold701/A _15044_/CLK _15044_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11207_ VGND VPWR VPWR VGND _11207_/X _11204_/X _11213_/S _11203_/X sky130_fd_sc_hd__mux2_1
X_12187_ VPWR VGND VGND VPWR _12187_/X hold291/A _12191_/B sky130_fd_sc_hd__or2_1
XFILLER_29_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11138_ VGND VPWR VGND VPWR _11138_/X _14890_/Q _11252_/A2 _11137_/X _11143_/S sky130_fd_sc_hd__o211a_1
X_13758__875 VPWR VGND VPWR VGND _15130_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_13951__1068 VPWR VGND VPWR VGND _15323_/CLK clkload26/A sky130_fd_sc_hd__inv_2
XFILLER_76_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11069_ VGND VPWR VGND VPWR _11069_/X _11068_/X _11067_/X _11176_/S _11185_/C1 sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_0_clk _12981__98/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_63_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13004__121 VPWR VGND VPWR VGND _14247_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_14828_ _14828_/Q _14832_/CLK _14828_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07300_ _07813_/A _15466_/Q _07300_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_14759_ hold287/A _14759_/CLK _14759_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08280_ VPWR VGND VPWR VGND _08277_/X _10061_/B _08280_/A2 _08280_/X _08280_/B2 sky130_fd_sc_hd__a22o_1
XFILLER_20_714 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07231_ VPWR VGND VGND VPWR _15445_/Q _08276_/B _08290_/B sky130_fd_sc_hd__nand2_1
X_07162_ VPWR VGND VGND VPWR _15473_/Q _07162_/B _07640_/A sky130_fd_sc_hd__nor2_1
X_07093_ VPWR VGND VPWR VGND _07372_/A _15451_/Q sky130_fd_sc_hd__inv_2
Xfanout204 VGND VPWR _12226_/A1 _12230_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout215 VGND VPWR fanout217/X _12256_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout237 VGND VPWR _12185_/A1 _12175_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09803_ VGND VPWR VPWR VGND _14249_/D fanout84/X _09830_/S hold377/X sky130_fd_sc_hd__mux2_1
Xfanout226 VGND VPWR _12863_/A1 _12720_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout248 VGND VPWR _12596_/C1 _12744_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_07995_ VGND VPWR VPWR VGND _15529_/D fanout34/X _08300_/S hold270/X sky130_fd_sc_hd__mux2_1
Xfanout259 VPWR VGND _12731_/S _12694_/S VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_55_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09734_ VGND VPWR VPWR VGND _14312_/D clone45/A _09757_/S hold262/X sky130_fd_sc_hd__mux2_1
XFILLER_39_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09665_ VGND VPWR VPWR VGND _14375_/D hold793/X _09687_/S fanout79/X sky130_fd_sc_hd__mux2_1
X_08616_ VGND VPWR VGND VPWR _15304_/D hold1054/X _08628_/A2 _08615_/X _11327_/A sky130_fd_sc_hd__o211a_1
X_09596_ VGND VPWR VPWR VGND _14472_/D clone49/A _09619_/S hold656/X sky130_fd_sc_hd__mux2_1
X_13551__668 VPWR VGND VPWR VGND _14882_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_08547_ VPWR VGND VGND VPWR _08554_/A _08554_/B _08548_/C sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_59_Left_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08478_ VPWR VGND VGND VPWR _08478_/X _15337_/Q _08482_/B sky130_fd_sc_hd__or2_1
X_07429_ VPWR VGND VGND VPWR _07429_/A _07539_/A _07429_/B sky130_fd_sc_hd__nand2_1
X_10440_ VGND VPWR VPWR VGND _10444_/B hold812/A _10554_/S hold696/A sky130_fd_sc_hd__mux2_1
XFILLER_7_718 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10371_ VGND VPWR VGND VPWR _10371_/X _10368_/X _10370_/X _10523_/A1 _10630_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_3_924 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12110_ VGND VPWR VGND VPWR _12110_/X _12109_/X _12108_/X _12118_/B1 _12115_/C1 sky130_fd_sc_hd__a211o_1
Xhold280 hold280/X hold280/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13445__562 VPWR VGND VPWR VGND _14720_/CLK clkload48/A sky130_fd_sc_hd__inv_2
X_12041_ VGND VPWR VGND VPWR _12041_/X _12038_/X _12040_/X _12226_/A1 _12202_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold291 hold291/X hold291/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout760 VPWR VGND _08002_/B1 _07426_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout793 VPWR VGND _08523_/B fanout802/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout782 VPWR VGND _07230_/S _07142_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout771 VGND VPWR _07418_/X _08104_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_1_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_58_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_73_474 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12874_ VGND VPWR VPWR VGND _15598_/D _07631_/X _14802_/D _15598_/Q sky130_fd_sc_hd__mux2_1
XANTENNA_120 _10893_/B1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_14613_ hold554/A _14613_/CLK _14613_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11825_ VPWR VGND VPWR VGND _11824_/X _12584_/A _12602_/B1 _11825_/X sky130_fd_sc_hd__a21o_1
X_15593_ _15593_/Q clkload49/A _15593_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_42_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14544_ hold586/A _14544_/CLK _14544_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11756_ VGND VPWR VPWR VGND _11756_/X hold586/A _11756_/S hold195/A sky130_fd_sc_hd__mux2_1
X_10707_ VPWR VGND VGND VPWR _10704_/X _10706_/X clone2/X _10707_/X sky130_fd_sc_hd__o21a_1
X_14475_ hold897/A _14475_/CLK _14475_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11687_ VGND VPWR VPWR VGND _11691_/B hold673/A _12052_/S hold253/A sky130_fd_sc_hd__mux2_1
X_10638_ VGND VPWR VPWR VGND _10642_/B hold515/A _10670_/S hold676/A sky130_fd_sc_hd__mux2_1
X_10569_ VGND VPWR VGND VPWR _10569_/X _10745_/A1 _10565_/X _10568_/X _10741_/C1 sky130_fd_sc_hd__o211a_1
X_12308_ VGND VPWR VPWR VGND _12312_/B hold720/A _12578_/S hold741/A sky130_fd_sc_hd__mux2_1
X_12239_ VGND VPWR VGND VPWR _12239_/X hold690/A _12705_/A2 _12256_/S _12238_/X sky130_fd_sc_hd__o211a_1
X_15027_ _15027_/Q _15027_/CLK _15027_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_69_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12950__67 VPWR VGND VPWR VGND _14193_/CLK clkload55/A sky130_fd_sc_hd__inv_2
XFILLER_39_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_29_1265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07780_ VPWR VGND VPWR VGND _08153_/B _07753_/B _07751_/X _08146_/B sky130_fd_sc_hd__a21o_1
XFILLER_49_460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xinput4 VGND VPWR input4/X ui_in[2] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_77_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09450_ VGND VPWR VGND VPWR _15581_/Q _09556_/C _15639_/Q _15580_/Q _09486_/C sky130_fd_sc_hd__and4bb_1
X_08401_ VGND VPWR VPWR VGND _15376_/D fanout10/X _08409_/S hold718/X sky130_fd_sc_hd__mux2_1
X_09381_ VPWR VGND VPWR VGND _09381_/X _09799_/A _09415_/B sky130_fd_sc_hd__or2_2
X_08332_ VGND VPWR VPWR VGND _15487_/D _09792_/A1 _08332_/S hold782/X sky130_fd_sc_hd__mux2_1
X_08263_ VPWR VGND VPWR VGND _08263_/A2 _07221_/X _08262_/X _08263_/X sky130_fd_sc_hd__a21o_1
X_07214_ VGND VPWR VGND VPWR _08201_/A _07369_/B _07369_/A sky130_fd_sc_hd__xnor2_4
X_13388__505 VPWR VGND VPWR VGND _14663_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_08194_ VPWR VGND VGND VPWR _08194_/B _08194_/Y _08690_/S sky130_fd_sc_hd__nand2_4
X_07145_ VPWR VGND VGND VPWR _14410_/Q _07304_/A2 _07304_/B1 _07145_/X sky130_fd_sc_hd__o21a_1
X_13429__546 VPWR VGND VPWR VGND _14704_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_10_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_43_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07978_ VGND VPWR VGND VPWR _15348_/Q clone13/X _15137_/Q _07978_/Y clone18/A sky130_fd_sc_hd__a22oi_4
X_09717_ VGND VPWR VPWR VGND _14326_/D fanout14/X _09728_/S hold739/X sky130_fd_sc_hd__mux2_1
X_13994__1111 VPWR VGND VPWR VGND _15366_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_14021__1138 VPWR VGND VPWR VGND _15393_/CLK clkload48/A sky130_fd_sc_hd__inv_2
X_09648_ VGND VPWR VPWR VGND _14422_/D hold1032/X _09659_/S fanout12/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1049 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12996__113 VPWR VGND VPWR VGND _14239_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
XFILLER_43_647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09579_ VGND VPWR VPWR VGND _14486_/D hold795/X _09590_/S fanout14/X sky130_fd_sc_hd__mux2_1
XFILLER_19_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12590_ VGND VPWR VPWR VGND _12590_/X _14374_/Q _12599_/S _14726_/Q sky130_fd_sc_hd__mux2_1
XFILLER_42_146 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11610_ VGND VPWR VGND VPWR _11610_/X _11638_/A1 _11606_/X _11609_/X _12115_/C1 sky130_fd_sc_hd__o211a_1
X_11541_ VPWR VGND _11542_/B _11541_/B _15431_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_13950__1067 VPWR VGND VPWR VGND _15322_/CLK clkload26/A sky130_fd_sc_hd__inv_2
XFILLER_51_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11472_ VGND VPWR VPWR VGND _11472_/X _15076_/Q _11475_/S _15074_/Q sky130_fd_sc_hd__mux2_1
X_14260_ hold730/A _14260_/CLK _14260_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14191_ _14191_/Q _14191_/CLK _14191_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10423_ VGND VPWR VGND VPWR _10423_/X _10667_/C1 _10418_/X _10422_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_10354_ VPWR VGND VGND VPWR _10354_/X _10685_/S _10354_/B sky130_fd_sc_hd__or2_1
XFILLER_65_1421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10285_ VPWR VGND VGND VPWR _10618_/A _10285_/B _10285_/Y sky130_fd_sc_hd__nor2_1
X_12024_ VPWR VGND VGND VPWR _12024_/X _12180_/S _12024_/B sky130_fd_sc_hd__or2_1
Xfanout590 VPWR VGND _09056_/S _09026_/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_59_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13222__339 VPWR VGND VPWR VGND _14497_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_34_614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12857_ VGND VPWR VPWR VGND _15581_/D _08072_/X _12877_/S _09240_/A sky130_fd_sc_hd__mux2_1
X_13573__690 VPWR VGND VPWR VGND _14904_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_11808_ VGND VPWR VPWR VGND _11808_/X hold962/A _12747_/S hold397/A sky130_fd_sc_hd__mux2_1
X_15576_ VGND VPWR VGND VPWR _15576_/Q _15576_/D clkload32/A sky130_fd_sc_hd__dfxtp_4
X_12788_ VGND VPWR VPWR VGND _12789_/B _08060_/B _12788_/S _08058_/B sky130_fd_sc_hd__mux2_1
X_14527_ hold228/A _14527_/CLK _14527_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13116__233 VPWR VGND VPWR VGND _14359_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_11739_ VGND VPWR VPWR VGND _11739_/X hold993/A _11748_/S hold556/A sky130_fd_sc_hd__mux2_1
X_14458_ hold566/A _14458_/CLK _14458_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14389_ _14389_/Q clkload22/A _14389_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_08950_ VPWR VGND VGND VPWR _08936_/X hold837/X _08933_/Y _15121_/Q hold838/A _11567_/A
+ sky130_fd_sc_hd__o221a_1
X_08881_ VGND VPWR VGND VPWR _15152_/D hold1239/X _08880_/B _08880_/Y _11308_/C1 sky130_fd_sc_hd__o211a_1
X_07901_ VGND VPWR VGND VPWR _07901_/X _07966_/A _10066_/B _07898_/Y _10071_/A sky130_fd_sc_hd__o211a_1
XFILLER_69_588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07832_ VGND VPWR _08155_/A _15549_/Q _15550_/Q _08208_/A VPWR VGND sky130_fd_sc_hd__and3_1
X_07763_ VPWR VGND VGND VPWR _15546_/Q _07773_/A _07772_/B sky130_fd_sc_hd__nand2_1
X_09502_ VGND VPWR VPWR VGND _14557_/D fanout40/X _09517_/S hold479/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13814__931 VPWR VGND VPWR VGND _15186_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XFILLER_77_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_912 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07694_ VGND VPWR _07694_/B _10066_/A _07694_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_77_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09433_ VGND VPWR VPWR VGND _14619_/D fanout32/X _09449_/S hold639/X sky130_fd_sc_hd__mux2_1
X_09364_ VGND VPWR VPWR VGND _14682_/D hold558/X _09379_/S fanout29/X sky130_fd_sc_hd__mux2_1
XFILLER_36_1022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08315_ VGND VPWR VPWR VGND _15504_/D fanout56/X _08318_/S hold1064/X sky130_fd_sc_hd__mux2_1
XANTENNA_31 _12829_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_20 _14389_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_09295_ VGND VPWR VPWR VGND _14746_/D fanout27/X _09302_/S hold193/X sky130_fd_sc_hd__mux2_1
XANTENNA_64 _09272_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_75 _09302_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08246_ VGND VPWR _15545_/Q _08246_/Y _15546_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
XANTENNA_53 _12869_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_42 _12866_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08177_ VPWR VGND VGND VPWR _08173_/Y _08176_/X _08017_/X _08214_/A _08177_/X _10058_/A1
+ sky130_fd_sc_hd__o221a_1
XANTENNA_86 _15468_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_97 fanout234/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07128_ VPWR VGND VPWR VGND _09198_/B _15639_/Q sky130_fd_sc_hd__inv_2
XFILLER_49_1438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10070_ VGND VPWR VPWR VGND _10071_/C _10069_/X _10068_/X _07654_/B _08287_/B _07410_/Y
+ sky130_fd_sc_hd__o2111a_1
XFILLER_43_1037 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_29_931 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13557__674 VPWR VGND VPWR VGND _14888_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_10972_ VGND VPWR VPWR VGND _10972_/X _14499_/Q _10972_/S hold480/A sky130_fd_sc_hd__mux2_1
X_12711_ VGND VPWR VGND VPWR _12711_/X _12708_/X _12710_/X _12748_/A1 _12744_/C1 sky130_fd_sc_hd__a211o_1
X_15430_ _15430_/Q clkload47/A _15430_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_989 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_31_617 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12642_ VGND VPWR VPWR VGND _12642_/X _14504_/Q _12651_/S _14184_/Q sky130_fd_sc_hd__mux2_1
XFILLER_24_680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12573_ VGND VPWR VPWR VGND _12573_/X _12570_/X _12581_/S _12569_/X sky130_fd_sc_hd__mux2_1
X_15361_ hold728/A _15361_/CLK _15361_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11524_ VGND VPWR VPWR VGND _11524_/X _11523_/X _11530_/S _15472_/Q sky130_fd_sc_hd__mux2_1
X_15292_ _15292_/Q _15292_/CLK _15292_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14312_ hold262/A _14312_/CLK _14312_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11455_ VGND VPWR VPWR VGND _11455_/X _11454_/X _11476_/S _15449_/Q sky130_fd_sc_hd__mux2_1
X_14243_ hold223/A _14243_/CLK _14243_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10406_ VPWR VGND VGND VPWR _10406_/X hold381/A _10702_/S sky130_fd_sc_hd__or2_1
XFILLER_7_378 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11386_ VGND VPWR VPWR VGND _11386_/X _14849_/Q _11392_/B _14817_/Q sky130_fd_sc_hd__mux2_1
X_14174_ _14174_/Q _14174_/CLK _14174_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10337_ VPWR VGND VGND VPWR _10334_/X _10336_/X _10765_/S _10337_/X sky130_fd_sc_hd__o21a_1
X_10268_ VGND VPWR VPWR VGND _10272_/B hold784/A _10609_/S hold449/A sky130_fd_sc_hd__mux2_1
XFILLER_79_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12920__37 VPWR VGND VPWR VGND _14163_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_12007_ VGND VPWR VGND VPWR _12007_/X _15010_/Q _12188_/A2 _11995_/S _12006_/X sky130_fd_sc_hd__o211a_1
XFILLER_79_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclone100 VGND VPWR _07890_/X clone100/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xclone111 VPWR VGND clone111/X _07659_/X VPWR VGND sky130_fd_sc_hd__buf_6
X_10199_ VGND VPWR VGND VPWR _10199_/X _11004_/A1 _10195_/X _10198_/X _11235_/C1 sky130_fd_sc_hd__o211a_1
Xclone133 VPWR VGND clone133/X fanout86/X VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_19_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15628_ _15628_/Q clkload49/A _15628_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15559_ _15559_/Q clkload43/A _15559_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08100_ VGND VPWR _08100_/B _12783_/B _08102_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_09080_ VGND VPWR VPWR VGND _15013_/D hold1107/X _09094_/S fanout25/X sky130_fd_sc_hd__mux2_1
X_13350__467 VPWR VGND VPWR VGND _14625_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_13993__1110 VPWR VGND VPWR VGND _15365_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_08031_ VPWR VGND VGND VPWR _08029_/X _08030_/X _08249_/B2 _08032_/C sky130_fd_sc_hd__o21a_1
X_14020__1137 VPWR VGND VPWR VGND _15392_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
Xhold802 hold802/X hold802/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/X hold846/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 hold835/X hold835/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold824 hold824/X hold824/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 hold813/X hold813/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 hold868/X hold868/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 hold879/X hold879/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ VGND VPWR _09986_/B _15607_/Q hold807/A _15608_/Q VPWR VGND sky130_fd_sc_hd__and3_1
Xhold857 hold857/X hold857/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ VPWR VGND VPWR VGND _08933_/Y _08933_/A sky130_fd_sc_hd__inv_2
XFILLER_44_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08864_ VPWR VGND VGND VPWR _08864_/X _15160_/Q _08868_/B sky130_fd_sc_hd__or2_1
X_13244__361 VPWR VGND VPWR VGND _14519_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_08795_ VGND VPWR VPWR VGND _15214_/D clone44/A _08808_/S hold172/X sky130_fd_sc_hd__mux2_1
X_07815_ VGND VPWR VPWR VGND _07820_/A _07815_/X _07815_/B sky130_fd_sc_hd__xor2_1
X_07746_ VGND VPWR _08096_/B _11535_/A _15553_/Q _07751_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_77_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_77_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07677_ VPWR VGND VPWR VGND _07676_/A _07119_/A clone17/X _07688_/A sky130_fd_sc_hd__a21oi_1
XFILLER_41_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09416_ VPWR VGND VPWR VGND _09416_/Y _09446_/S sky130_fd_sc_hd__inv_2
XFILLER_41_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_55_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_32_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09347_ VPWR VGND VGND VPWR hold1372/X _09357_/S _09347_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_8_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09278_ VPWR VGND VGND VPWR _09278_/X _09278_/A _09307_/S sky130_fd_sc_hd__or2_1
X_08229_ VPWR VGND VPWR VGND _08228_/X _08214_/X _08217_/X _08230_/B _08294_/B1 sky130_fd_sc_hd__a22o_1
XFILLER_10_1014 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11240_ VGND VPWR VPWR VGND _11240_/X _14218_/Q _11240_/S _15226_/Q sky130_fd_sc_hd__mux2_1
X_11171_ VPWR VGND VPWR VGND _11170_/X _11181_/A1 _11169_/X _11171_/Y sky130_fd_sc_hd__a21oi_1
X_10122_ VGND VPWR VPWR VGND _10122_/X hold780/A _10353_/S hold318/A sky130_fd_sc_hd__mux2_1
XFILLER_76_845 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14930_ _14930_/Q clkload29/A _14930_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10053_ VPWR VGND VGND VPWR _14803_/Q _10053_/Y _10053_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14861_ _15701_/A clkload25/A _14861_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1395 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14792_ hold661/A _14792_/CLK _14792_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_73_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10955_ VPWR VGND VGND VPWR _10955_/X hold834/A _11142_/S sky130_fd_sc_hd__or2_1
X_10886_ VGND VPWR VPWR VGND _10886_/X _15387_/Q _11109_/S _15534_/Q sky130_fd_sc_hd__mux2_1
X_15413_ hold375/A _15413_/CLK _15413_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12625_ VPWR VGND VGND VPWR _12625_/X hold540/A _12635_/B sky130_fd_sc_hd__or2_1
X_15344_ _15344_/Q _15344_/CLK _15344_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_40_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12556_ VGND VPWR VPWR VGND _12556_/X hold737/A _12671_/S hold385/A sky130_fd_sc_hd__mux2_1
X_11507_ VGND VPWR VPWR VGND _15086_/D _11506_/X _11538_/S hold1427/X sky130_fd_sc_hd__mux2_1
X_13187__304 VPWR VGND VPWR VGND _14462_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_15275_ hold895/A _15275_/CLK _15275_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12487_ VPWR VGND VGND VPWR _12487_/X hold301/A _12716_/S sky130_fd_sc_hd__or2_1
X_11438_ VGND VPWR VGND VPWR _11438_/X _14934_/Q _11303_/A _11439_/A2 sky130_fd_sc_hd__a21bo_1
X_14226_ hold213/A _14226_/CLK _14226_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14157_ hold636/A _14157_/CLK _14157_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11369_ VGND VPWR VPWR VGND _11369_/X _11364_/X _11387_/S _14844_/Q sky130_fd_sc_hd__mux2_1
X_13228__345 VPWR VGND VPWR VGND _14503_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
XFILLER_26_1032 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08580_ VGND VPWR _08580_/B _08580_/Y _08580_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07600_ VPWR VGND VPWR VGND _15637_/Q _07929_/A2 _07600_/X _07908_/B1 _07519_/B _07599_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_78_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07531_ VGND VPWR _07531_/X _07531_/B _07531_/A _07531_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_74_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07462_ VPWR VGND VGND VPWR _07462_/A _08603_/A _07462_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_1448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09201_ VGND VPWR VPWR VGND _14892_/D hold1073/X _09213_/S clone133/X sky130_fd_sc_hd__mux2_1
X_07393_ _07306_/B _15465_/Q _07878_/A _07876_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_09132_ _14966_/D fanout91/X fanout87/X _09130_/Y _09131_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09063_ _15030_/D fanout93/X fanout89/X _09090_/S _09062_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08014_ VGND VPWR VGND VPWR _08013_/X _08014_/X _08014_/A _08014_/B sky130_fd_sc_hd__or3b_4
Xhold621 hold621/X hold621/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold610 hold610/X hold610/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold632 hold632/X hold632/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 hold654/X hold654/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 hold643/X hold643/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 hold665/X hold665/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 hold676/X hold676/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 hold687/X hold687/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 hold698/X hold698/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ VPWR VGND VPWR VGND _09965_/X _15571_/Q _12846_/B sky130_fd_sc_hd__or2_2
X_09896_ VPWR VGND VPWR VGND _09895_/X _08857_/Y _09893_/Y _14145_/D hold149/X sky130_fd_sc_hd__a22o_1
X_08916_ VPWR VGND VGND VPWR _08916_/X _15134_/Q _08926_/B sky130_fd_sc_hd__or2_1
Xhold1343 _09998_/B _09997_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 _10016_/A _15622_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 hold1332/X _15085_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1310 _09981_/B _15607_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08847_ VGND VPWR VPWR VGND _15166_/D _09228_/A0 _08847_/S hold842/X sky130_fd_sc_hd__mux2_1
Xhold1376 _07601_/A _15544_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1354 hold1354/X _15299_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1365 hold1365/X _14666_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1387 hold1387/X _15152_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1398 hold1398/X _15353_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_40_Left_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08778_ VGND VPWR VPWR VGND _15228_/D fanout98/X _08779_/S hold318/X sky130_fd_sc_hd__mux2_1
X_07729_ VPWR VGND VPWR VGND _07827_/D _15585_/Q _07714_/X _07730_/B sky130_fd_sc_hd__a21o_1
X_13021__138 VPWR VGND VPWR VGND _14264_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
XFILLER_25_263 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10740_ VGND VPWR VGND VPWR _10740_/X hold926/A _10744_/A2 _10739_/X _10588_/S sky130_fd_sc_hd__o211a_1
X_10671_ VGND VPWR VGND VPWR _10671_/X _10670_/X _10669_/X _10557_/A _10717_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_16_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_16_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12410_ VGND VPWR VGND VPWR _12410_/X _15503_/Q _12743_/A2 _12721_/S _12409_/X sky130_fd_sc_hd__o211a_1
X_13669__786 VPWR VGND VPWR VGND _15009_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_12341_ VGND VPWR VGND VPWR _12341_/X _12338_/X _12340_/X _12588_/A1 _12744_/C1 sky130_fd_sc_hd__a211o_1
Xclone54 VGND VPWR clone54/X clone55/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_12272_ VGND VPWR VPWR VGND _12272_/X _14494_/Q _12282_/S _14174_/Q sky130_fd_sc_hd__mux2_1
X_15060_ hold624/A _15060_/CLK _15060_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11223_ VGND VPWR VPWR VGND _11223_/X hold841/A _11223_/S hold509/A sky130_fd_sc_hd__mux2_1
XFILLER_4_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11154_ VPWR VGND VPWR VGND _11153_/X _11247_/A _12713_/B1 _11154_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11085_ VPWR VGND VGND VPWR _11085_/X _15254_/Q _11091_/S sky130_fd_sc_hd__or2_1
XFILLER_27_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10105_ VGND VPWR VGND VPWR _10105_/X hold922/A _10629_/A2 _10104_/X _10614_/A1 sky130_fd_sc_hd__o211a_1
X_14913_ hold585/A _14913_/CLK _14913_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10036_ VPWR VGND VGND VPWR _10038_/C _10036_/B _15630_/D sky130_fd_sc_hd__nor2_1
XFILLER_7_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_75_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14844_ _14844_/Q clkload19/A _14844_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14775_ hold485/A _14775_/CLK _14775_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11987_ VPWR VGND VGND VPWR _11987_/X _11995_/S _11987_/B sky130_fd_sc_hd__or2_1
X_13613__730 VPWR VGND VPWR VGND _14953_/CLK clkload53/A sky130_fd_sc_hd__inv_2
XFILLER_44_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10938_ VPWR VGND VGND VPWR _10938_/X _11170_/S _10938_/B sky130_fd_sc_hd__or2_1
XFILLER_32_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_907 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10869_ VGND VPWR VPWR VGND _10869_/X _14464_/Q _10885_/S _14752_/Q sky130_fd_sc_hd__mux2_1
XFILLER_31_299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12608_ VPWR VGND VGND VPWR _12608_/X _12624_/S _12608_/B sky130_fd_sc_hd__or2_1
X_15327_ _15327_/Q _15327_/CLK _15327_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14195__913 _14195_/D _14195__913/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_12539_ VGND VPWR VPWR VGND _12539_/X hold575/A _12539_/S hold373/A sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15258_ _15258_/Q _15258_/CLK _15258_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14209_ _14209_/Q _14209_/CLK _14209_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15189_ hold737/A _15189_/CLK _15189_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13462__579 VPWR VGND VPWR VGND _14737_/CLK clkload55/A sky130_fd_sc_hd__inv_2
Xfanout419 VGND VPWR fanout424/X _11254_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout408 VGND VPWR _10622_/C1 _10630_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09750_ VGND VPWR VPWR VGND _14296_/D fanout19/X _09756_/S hold514/X sky130_fd_sc_hd__mux2_1
X_08701_ VGND VPWR VGND VPWR _15281_/D hold1059/X _08701_/A2 _08700_/X _11937_/C1
+ sky130_fd_sc_hd__o211a_1
X_09681_ VGND VPWR VPWR VGND _14359_/D hold1038/X _09693_/S fanout17/X sky130_fd_sc_hd__mux2_1
X_08632_ VPWR VGND VPWR VGND _15298_/Q _08700_/A2 _08632_/X _08711_/B1 _08631_/X _08700_/B1
+ sky130_fd_sc_hd__a221o_1
XFILLER_78_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08563_ VGND VPWR VGND VPWR _08563_/X _08605_/A _08615_/B1 hold886/X _08562_/Y sky130_fd_sc_hd__a211o_1
XFILLER_35_550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08494_ VGND VPWR VGND VPWR _08495_/A2 _15638_/Q _09937_/B _08493_/Y sky130_fd_sc_hd__a21oi_2
X_07514_ VPWR VGND _07515_/A _07519_/B _15466_/Q VPWR VGND sky130_fd_sc_hd__xor2_2
X_13356__473 VPWR VGND VPWR VGND _14631_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
XFILLER_22_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07445_ VPWR VGND VGND VPWR _07447_/A _15456_/Q _07714_/A sky130_fd_sc_hd__or2_1
Xfanout15 VGND VPWR _08070_/X fanout15/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout37 VGND VPWR _07976_/X fanout37/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout26 VGND VPWR fanout26/X _08032_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout48 VPWR VGND VGND VPWR _07890_/X fanout48/X sky130_fd_sc_hd__buf_8
XFILLER_52_1423 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_918 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07376_ VPWR VGND VGND VPWR _07376_/A _07376_/B _07376_/Y sky130_fd_sc_hd__nor2_1
X_09115_ VGND VPWR VPWR VGND _14980_/D hold335/X _09125_/S fanout21/X sky130_fd_sc_hd__mux2_1
X_12956__73 VPWR VGND VPWR VGND _14199_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_09046_ VGND VPWR VPWR VGND _15044_/D hold701/X _09056_/S _08051_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold462 hold462/X hold462/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1186 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold440 hold440/X hold440/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 hold451/X hold451/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/X hold495/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 hold484/X hold484/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold473/X hold473/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09948_ VGND VPWR _09947_/C _14128_/Q _09949_/B _14129_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
X_09879_ VPWR VGND VPWR VGND _09878_/Y _09877_/X _09882_/A _14150_/D sky130_fd_sc_hd__a21oi_1
Xhold1140 hold1140/X _14241_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 hold1151/X _14593_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _14148_/D _09884_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 hold1162/X _15341_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1184 hold1184/X _14689_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ VGND VPWR VPWR VGND _11910_/X hold730/A _12227_/S hold292/A sky130_fd_sc_hd__mux2_1
Xhold1195 hold1195/X _14630_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ VGND VPWR VPWR VGND _11841_/X _11838_/X _12100_/S _11837_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14560_ _14560_/Q _14560_/CLK _14560_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_54_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11772_ VGND VPWR VPWR VGND _11772_/X hold779/A _12155_/S hold494/A sky130_fd_sc_hd__mux2_1
XFILLER_14_723 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_41_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10723_ VGND VPWR VPWR VGND _10723_/X hold617/A _10743_/B hold211/A sky130_fd_sc_hd__mux2_1
X_14491_ _14491_/Q _14491_/CLK _14491_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10654_ VGND VPWR VPWR VGND _10655_/B _10653_/Y clone2/A _10645_/Y sky130_fd_sc_hd__mux2_1
XFILLER_13_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10585_ VGND VPWR VGND VPWR _10585_/X _10584_/X _10583_/X _10745_/A1 _10741_/C1 sky130_fd_sc_hd__a211o_1
Xclkload29 VGND VPWR VGND VPWR clkload29/Y clkload29/A sky130_fd_sc_hd__inv_8
X_15112_ hold758/A _15112_/CLK _15112_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12324_ VGND VPWR VPWR VGND _12325_/B _12323_/Y _12583_/S _12315_/Y sky130_fd_sc_hd__mux2_1
Xclkload18 VGND VPWR VPWR VGND clkload18/A clkload18/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_68_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12255_ VGND VPWR VGND VPWR _12255_/X _12581_/S _12252_/X _12254_/X _12572_/C1 sky130_fd_sc_hd__o211a_1
X_15043_ hold402/A _15043_/CLK _15043_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11206_ VGND VPWR VGND VPWR _11206_/X _11215_/C1 _11202_/X _11205_/X _11217_/C1 sky130_fd_sc_hd__o211a_1
X_12186_ VGND VPWR VPWR VGND _12186_/X hold528/A _12191_/B hold270/A sky130_fd_sc_hd__mux2_1
X_11137_ VPWR VGND VGND VPWR _11137_/X hold363/A _11146_/B sky130_fd_sc_hd__or2_1
XFILLER_77_940 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13299__416 VPWR VGND VPWR VGND _14574_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
XFILLER_76_450 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11068_ VGND VPWR VPWR VGND _11068_/X hold935/A _11068_/S hold310/A sky130_fd_sc_hd__mux2_1
XFILLER_64_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_697 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10019_ VPWR VGND VGND VPWR _10021_/B _10019_/B _15623_/D sky130_fd_sc_hd__nor2_1
X_13043__160 VPWR VGND VPWR VGND _14286_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_14827_ _14827_/Q _14832_/CLK _14827_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14758_ _14758_/Q _14758_/CLK _14758_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_36_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14689_ _14689_/Q _14689_/CLK _14689_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07230_ VGND VPWR VPWR VGND _07230_/S _15590_/Q _14379_/Q _08290_/B sky130_fd_sc_hd__mux2_2
X_07161_ VPWR VGND _07163_/A _07162_/B _15473_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07092_ VPWR VGND VPWR VGND _07371_/A _15452_/Q sky130_fd_sc_hd__inv_2
Xfanout205 VGND VPWR _07978_/Y _12226_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout238 VPWR VGND _12185_/A1 _12193_/C1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout227 VPWR VGND _12863_/A1 fanout234/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout216 VGND VPWR fanout217/X _12580_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09802_ _14250_/D fanout91/X fanout87/X _09800_/Y _09801_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xfanout249 VGND VPWR _12596_/C1 _12703_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_07994_ VGND VPWR VGND VPWR _07994_/X _07991_/X _07994_/C _07994_/B _07994_/A sky130_fd_sc_hd__or4b_4
XFILLER_45_1260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13919__1036 VPWR VGND VPWR VGND _15291_/CLK clkload16/A sky130_fd_sc_hd__inv_2
XFILLER_80_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09733_ VGND VPWR VPWR VGND _14313_/D fanout85/X _09760_/S hold323/X sky130_fd_sc_hd__mux2_1
XFILLER_41_1168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09664_ VGND VPWR VPWR VGND _09687_/S hold1194/X clone49/X _14376_/D sky130_fd_sc_hd__mux2_2
X_08615_ VGND VPWR VGND VPWR _08615_/X _08617_/A _08615_/B1 hold986/X _08614_/Y sky130_fd_sc_hd__a211o_1
X_09595_ VGND VPWR VPWR VGND _14473_/D fanout85/X _09619_/S hold604/X sky130_fd_sc_hd__mux2_1
X_08546_ VPWR VGND _08554_/B _08546_/B _08546_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08477_ VGND VPWR VGND VPWR _15338_/D hold1137/X _08483_/A2 _08476_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_13092__209 VPWR VGND VPWR VGND _14335_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_07428_ VPWR VGND VGND VPWR _07429_/B _15467_/Q _07519_/B sky130_fd_sc_hd__or2_1
X_07359_ VPWR VGND VPWR VGND _08180_/A _08223_/A _08201_/A _08162_/A _10061_/C sky130_fd_sc_hd__or4_1
X_10370_ VGND VPWR VGND VPWR _10370_/X _15488_/Q _10633_/A2 _10369_/X _10625_/S sky130_fd_sc_hd__o211a_1
X_09029_ VGND VPWR VPWR VGND _15061_/D hold509/X _09053_/S fanout83/X sky130_fd_sc_hd__mux2_1
Xhold270 hold270/X hold270/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ VGND VPWR VGND VPWR _12040_/X hold844/A _12040_/A2 _11925_/S _12039_/X sky130_fd_sc_hd__o211a_1
Xhold281 hold281/X hold281/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/X hold292/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13790__907 VPWR VGND VPWR VGND _15162_/CLK clkload25/A sky130_fd_sc_hd__inv_2
Xfanout750 VPWR VGND _07552_/B1 _07534_/Y VPWR VGND sky130_fd_sc_hd__buf_2
X_13027__144 VPWR VGND VPWR VGND _14270_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
Xfanout761 VPWR VGND _08299_/A2 _08249_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout783 VGND VPWR _07142_/X _07220_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout772 VGND VPWR _08066_/B _10075_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout794 VPWR VGND _08714_/A2 _08667_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
X_13831__948 VPWR VGND VPWR VGND _15203_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
XFILLER_45_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12873_ VGND VPWR VPWR VGND _15597_/D _07645_/X _14802_/D _15597_/Q sky130_fd_sc_hd__mux2_1
XANTENNA_110 _10737_/C1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_14612_ hold677/A _14612_/CLK _14612_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_121 _10893_/B1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11824_ VPWR VGND _11824_/X _11823_/X _11819_/X _12583_/S _11815_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15592_ _15592_/Q clkload49/A _15592_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14543_ hold804/A _14543_/CLK _14543_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11755_ VGND VPWR VPWR VGND _11755_/X hold689/A _12086_/S hold221/A sky130_fd_sc_hd__mux2_1
X_10706_ VGND VPWR VGND VPWR _10706_/X _10703_/A _10702_/X _10705_/X _10706_/C1 sky130_fd_sc_hd__o211a_1
X_13684__801 VPWR VGND VPWR VGND _15024_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_14474_ _14474_/Q _14474_/CLK _14474_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11686_ VPWR VGND VPWR VGND _11685_/X _12722_/A1 _11684_/X _11686_/Y sky130_fd_sc_hd__a21oi_1
X_10637_ VPWR VGND VGND VPWR _10618_/Y _10636_/X _10710_/B _14393_/Q _14393_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
X_13725__842 VPWR VGND VPWR VGND _15097_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_10568_ VPWR VGND VGND VPWR _10568_/X _10588_/S _10568_/B sky130_fd_sc_hd__or2_1
X_12307_ VPWR VGND VGND VPWR _12288_/Y _12306_/X _12269_/B _15464_/Q _15464_/D _11341_/A
+ sky130_fd_sc_hd__o221a_1
X_10499_ VGND VPWR VPWR VGND _10499_/X hold459/A _10516_/S hold410/A sky130_fd_sc_hd__mux2_1
X_15026_ _15026_/Q _15026_/CLK _15026_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12238_ VPWR VGND VGND VPWR _12238_/X hold182/A _12318_/S sky130_fd_sc_hd__or2_1
X_12169_ VGND VPWR VPWR VGND _12169_/X hold943/A _12171_/S hold196/A sky130_fd_sc_hd__mux2_1
XFILLER_49_472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08400_ VGND VPWR VPWR VGND _15377_/D fanout13/X _08411_/S hold802/X sky130_fd_sc_hd__mux2_1
XFILLER_75_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09380_ VPWR VGND VGND VPWR _09415_/B _15580_/Q _09556_/C _09240_/A sky130_fd_sc_hd__nand3b_1
XFILLER_51_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08331_ VGND VPWR VPWR VGND _15488_/D _09548_/A1 _08338_/S hold1061/X sky130_fd_sc_hd__mux2_1
XFILLER_60_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08262_ VPWR VGND VPWR VGND _10061_/A _08280_/A2 _08262_/X _08293_/B1 _15067_/Q _08261_/X
+ sky130_fd_sc_hd__a221o_1
X_07213_ VPWR VGND _07213_/X _07369_/B _15450_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_08193_ VPWR VGND VPWR VGND _08252_/A2 _15158_/Q _08192_/X _08193_/X sky130_fd_sc_hd__a21o_1
X_07144_ VPWR VGND VPWR VGND _07144_/A1 _08294_/B1 _07144_/X wire858/X _15576_/Q _07714_/A
+ sky130_fd_sc_hd__a221o_1
X_13468__585 VPWR VGND VPWR VGND _14743_/CLK clkload9/A sky130_fd_sc_hd__inv_2
XFILLER_10_15 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12926__43 VPWR VGND VPWR VGND _14169_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_07977_ VGND VPWR VPWR VGND _15530_/D fanout37/X _08267_/S hold266/X sky130_fd_sc_hd__mux2_1
X_09716_ VGND VPWR VPWR VGND _14327_/D fanout15/X _09728_/S hold850/X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_55_442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09647_ VGND VPWR VPWR VGND _14423_/D hold887/X _09659_/S fanout15/X sky130_fd_sc_hd__mux2_1
X_09578_ VGND VPWR VPWR VGND _14487_/D hold763/X _09590_/S fanout16/X sky130_fd_sc_hd__mux2_1
X_08529_ VPWR VGND _15322_/D _08529_/B _08529_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_35_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_19_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11540_ VPWR VGND VPWR VGND _11539_/Y _11541_/B _11542_/A _15430_/D sky130_fd_sc_hd__a21oi_1
XFILLER_19_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13709__826 VPWR VGND VPWR VGND _15049_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_11471_ VGND VPWR VPWR VGND _15074_/D _11470_/X _11477_/S _15074_/Q sky130_fd_sc_hd__mux2_1
X_14190_ _14190_/Q _14190_/CLK _14190_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10422_ VGND VPWR VGND VPWR _10422_/X _10421_/X _10420_/X _10652_/S _10717_/C1 sky130_fd_sc_hd__a211o_1
X_10353_ VGND VPWR VPWR VGND _10353_/X _14450_/Q _10353_/S hold282/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12023_ VGND VPWR VPWR VGND _12023_/X _14455_/Q _12190_/S hold659/A sky130_fd_sc_hd__mux2_1
X_10284_ VGND VPWR VPWR VGND _10285_/B _10283_/Y _10617_/S _10275_/Y sky130_fd_sc_hd__mux2_1
XFILLER_66_718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout580 _09269_/S _09272_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_59_792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout591 VPWR VGND _08850_/S _08842_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_13261__378 VPWR VGND VPWR VGND _14536_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_12856_ VGND VPWR VPWR VGND _15580_/D _08093_/X _12877_/S _09311_/B sky130_fd_sc_hd__mux2_1
X_11807_ VPWR VGND VGND VPWR _12584_/A _11807_/B _11807_/Y sky130_fd_sc_hd__nor2_1
X_15575_ _15575_/Q clkload43/A _15575_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_873 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12787_ VPWR VGND VPWR VGND _12878_/C _08571_/Y _12786_/X _15554_/D sky130_fd_sc_hd__a21oi_1
X_14526_ hold209/A _14526_/CLK _14526_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13155__272 VPWR VGND VPWR VGND _14430_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_13918__1035 VPWR VGND VPWR VGND _15290_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_11738_ VGND VPWR VGND VPWR _11738_/X hold832/A _12488_/A2 _12720_/A1 _11737_/X sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_78_Left_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11669_ VPWR VGND VGND VPWR _11669_/X hold188/A _11965_/S sky130_fd_sc_hd__or2_1
X_14457_ _14457_/Q _14457_/CLK _14457_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14388_ _14388_/Q clkload17/A _14388_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_51_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08880_ VPWR VGND VGND VPWR _08880_/A _08880_/Y _08880_/B sky130_fd_sc_hd__nand2_1
X_15009_ _15009_/Q _15009_/CLK _15009_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07900_ VPWR VGND _10066_/B _07900_/B _07900_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_13502__619 VPWR VGND VPWR VGND _14777_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_07831_ VPWR VGND _08208_/A _08220_/B _15548_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_57_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07762_ VPWR VGND VPWR VGND _07826_/D _15593_/Q _07765_/B _07772_/B _09311_/B sky130_fd_sc_hd__a22o_1
X_09501_ VGND VPWR VPWR VGND _14558_/D clone6/X _09514_/S hold490/X sky130_fd_sc_hd__mux2_1
X_13853__970 VPWR VGND VPWR VGND _15225_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_77_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07693_ VGND VPWR _07693_/B _07693_/Y _07693_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_37_486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09432_ VGND VPWR VPWR VGND _14620_/D fanout36/X _09441_/S hold618/X sky130_fd_sc_hd__mux2_1
X_09363_ VGND VPWR VPWR VGND _14683_/D hold536/X _09377_/S fanout33/X sky130_fd_sc_hd__mux2_1
XFILLER_21_821 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08314_ VGND VPWR VPWR VGND _15505_/D fanout63/X _08335_/S hold1060/X sky130_fd_sc_hd__mux2_1
XANTENNA_32 _08730_/B1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_21 _14389_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_09294_ VGND VPWR VPWR VGND _14747_/D fanout31/X _09310_/S hold242/X sky130_fd_sc_hd__mux2_1
XANTENNA_10 _08212_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_43 fanout282/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_65 _09272_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08245_ VGND VPWR VGND VPWR _08245_/X _08280_/A2 _08242_/X _10062_/A _08244_/X sky130_fd_sc_hd__a211o_1
XFILLER_36_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_54 _11209_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08176_ VPWR VGND VPWR VGND clone20/A _15159_/Q _08175_/X _08176_/X sky130_fd_sc_hd__a21o_1
XANTENNA_76 _09091_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_87 _15474_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_98 fanout234/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07127_ VPWR VGND VPWR VGND _15606_/D hold807/X sky130_fd_sc_hd__inv_2
XFILLER_48_718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13098__215 VPWR VGND VPWR VGND _14341_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_10971_ VGND VPWR VPWR VGND _10975_/B hold623/A _10972_/S hold400/A sky130_fd_sc_hd__mux2_1
XFILLER_71_732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_46_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12710_ VGND VPWR VGND VPWR _12710_/X _15029_/Q _12746_/A2 _11810_/S _12709_/X sky130_fd_sc_hd__o211a_1
XFILLER_15_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12641_ VGND VPWR VPWR VGND _12645_/B _14632_/Q _12661_/S _14664_/Q sky130_fd_sc_hd__mux2_1
X_13139__256 VPWR VGND VPWR VGND _14414_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_12572_ VGND VPWR VGND VPWR _12572_/X _12580_/A1 _12568_/X _12571_/X _12572_/C1 sky130_fd_sc_hd__o211a_1
X_15360_ _15360_/Q _15360_/CLK _15360_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11523_ VGND VPWR VPWR VGND _11523_/X _15093_/Q _11529_/S _15091_/Q sky130_fd_sc_hd__mux2_1
X_15291_ _15291_/Q _15291_/CLK _15291_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14311_ _14311_/Q _14311_/CLK _14311_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11454_ VGND VPWR VPWR VGND _11454_/X _15070_/Q _11490_/S _15068_/Q sky130_fd_sc_hd__mux2_1
XFILLER_7_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14242_ hold198/A _14242_/CLK _14242_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10405_ VGND VPWR VPWR VGND _10405_/X hold680/A _10702_/S hold271/A sky130_fd_sc_hd__mux2_1
X_14173_ hold855/A _14173_/CLK _14173_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11385_ VGND VPWR VPWR VGND _14848_/D _11384_/X _11388_/S hold1300/X sky130_fd_sc_hd__mux2_1
X_10336_ VGND VPWR VGND VPWR _10336_/X _11110_/A _10332_/X _10335_/X _11096_/C1 sky130_fd_sc_hd__o211a_1
X_13796__913 VPWR VGND VPWR VGND _15168_/CLK clkload13/A sky130_fd_sc_hd__inv_2
XFILLER_3_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10267_ VPWR VGND VGND VPWR _10248_/Y _10266_/X _12380_/B _14383_/Q _14383_/D _12492_/C1
+ sky130_fd_sc_hd__o221a_1
X_12006_ VPWR VGND VGND VPWR _12006_/X hold343/A _12006_/B sky130_fd_sc_hd__or2_1
XFILLER_39_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10198_ VPWR VGND VGND VPWR _10198_/X _10995_/S _10198_/B sky130_fd_sc_hd__or2_1
X_13837__954 VPWR VGND VPWR VGND _15209_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_47_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_46_261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15627_ _15627_/Q clkload49/A _15627_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_979 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12839_ VGND VPWR _15567_/Q _15569_/Q _12840_/B _15568_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_21_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15558_ _15558_/Q clkload44/A _15558_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14509_ hold188/A _14509_/CLK _14509_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15489_ hold821/A _15489_/CLK _15489_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08030_ VPWR VGND VPWR VGND _08027_/X _08025_/A _07414_/Y _08030_/X _08280_/B2 sky130_fd_sc_hd__a22o_1
Xhold803 hold803/X hold803/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 hold814/X hold814/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 hold825/X hold825/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 hold836/X hold836/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 hold847/X hold847/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 hold869/X hold869/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ VGND VPWR VPWR VGND hold807/A _09981_/X _09981_/B sky130_fd_sc_hd__xor2_1
Xhold858 hold858/X hold858/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08932_ VPWR VGND _08932_/X _09892_/A _08935_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08863_ VGND VPWR VPWR VGND _09893_/A _08862_/C _09970_/A _08863_/X sky130_fd_sc_hd__or3b_1
XFILLER_57_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08794_ VGND VPWR VPWR VGND _15215_/D fanout47/X _08808_/S hold274/X sky130_fd_sc_hd__mux2_1
X_07814_ _07815_/B _07859_/A _07813_/A _07813_/B _07296_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07745_ VPWR VGND VPWR VGND _07751_/C _11535_/A _15553_/Q _07745_/X sky130_fd_sc_hd__a21o_1
XFILLER_77_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09415_ VPWR VGND VGND VPWR _09415_/B _09415_/Y _09694_/A sky130_fd_sc_hd__nor2_2
X_07676_ VPWR VGND VPWR VGND _07676_/Y _07676_/A sky130_fd_sc_hd__inv_2
XFILLER_53_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13630__747 VPWR VGND VPWR VGND _14970_/CLK clkload37/A sky130_fd_sc_hd__inv_2
XFILLER_12_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09346_ VGND VPWR VGND VPWR _09660_/B _09799_/A _09346_/X sky130_fd_sc_hd__or2_4
X_09277_ VPWR VGND VPWR VGND _09277_/Y _09307_/S sky130_fd_sc_hd__inv_2
X_08228_ VGND VPWR VGND VPWR _08228_/X _08280_/A2 _08225_/X _08223_/A _08227_/X sky130_fd_sc_hd__a211o_1
X_13483__600 VPWR VGND VPWR VGND _14758_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_08159_ VPWR VGND VGND VPWR _08180_/C _08201_/A _08201_/C sky130_fd_sc_hd__or2_1
X_11170_ VGND VPWR VPWR VGND _11170_/X _11167_/X _11170_/S _11166_/X sky130_fd_sc_hd__mux2_1
X_13524__641 VPWR VGND VPWR VGND _14799_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_10121_ VGND VPWR VPWR VGND _10121_/X _14476_/Q _10612_/S hold396/A sky130_fd_sc_hd__mux2_1
X_10052_ VGND VPWR VGND VPWR _14803_/Q _11117_/B _10053_/B sky130_fd_sc_hd__and2_4
X_13917__1034 VPWR VGND VPWR VGND _15289_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_14860_ _15702_/A clkload26/A _14860_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1330 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_29_751 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14791_ hold670/A _14791_/CLK _14791_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_21_1177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10954_ VGND VPWR VPWR VGND _10954_/X _10953_/X _11170_/S _10952_/X sky130_fd_sc_hd__mux2_1
X_10885_ VGND VPWR VPWR VGND _10885_/X _15020_/Q _10885_/S hold748/A sky130_fd_sc_hd__mux2_1
X_12624_ VGND VPWR VPWR VGND _12624_/X _12623_/X _12624_/S _12622_/X sky130_fd_sc_hd__mux2_1
X_15412_ hold488/A _15412_/CLK _15412_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15343_ _15343_/Q _15343_/CLK _15343_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12555_ VGND VPWR VGND VPWR _12555_/X _12656_/A1 _12554_/X _12551_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_11506_ VGND VPWR VPWR VGND _11506_/X _11505_/X _11537_/S _15466_/Q sky130_fd_sc_hd__mux2_1
XFILLER_12_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15274_ hold915/A _15274_/CLK _15274_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12486_ VGND VPWR VPWR VGND _12486_/X hold416/A _12716_/S hold542/A sky130_fd_sc_hd__mux2_1
X_11437_ VGND VPWR VGND VPWR _14933_/D hold1345/X _11439_/A2 _11436_/X _11347_/A sky130_fd_sc_hd__o211a_1
X_14225_ hold308/A _14225_/CLK _14225_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11368_ VGND VPWR VGND VPWR _11387_/S _11356_/X _11368_/C _11368_/B _11368_/A sky130_fd_sc_hd__or4b_4
X_14156_ hold396/A _14156_/CLK _14156_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10319_ VGND VPWR VGND VPWR _10319_/X _10316_/X _10318_/X _11112_/A _11263_/C1 sky130_fd_sc_hd__a211o_1
X_13267__384 VPWR VGND VPWR VGND _14542_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_11299_ VGND VPWR VPWR VGND _11300_/B _14818_/Q _11299_/S _14386_/Q sky130_fd_sc_hd__mux2_1
XFILLER_67_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_1127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_43_1391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_78_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07530_ VPWR VGND VPWR VGND _07530_/B _07530_/C _07530_/A _07531_/A sky130_fd_sc_hd__or3_4
X_14989_ hold589/A _14989_/CLK _14989_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_74_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07461_ VPWR VGND VGND VPWR _07462_/B _15451_/Q _15596_/Q sky130_fd_sc_hd__or2_1
XFILLER_35_776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07392_ VPWR VGND VGND VPWR _07297_/B _15467_/Q _07819_/A sky130_fd_sc_hd__nand2b_1
X_09200_ _14893_/D fanout91/X fanout87/X _09213_/S _09199_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_37_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09131_ VPWR VGND VGND VPWR _09131_/X _09131_/A _09157_/S sky130_fd_sc_hd__or2_1
X_09062_ VPWR VGND VGND VPWR hold1410/X _09090_/S _09062_/Y sky130_fd_sc_hd__nand2b_1
X_08013_ VPWR VGND _08013_/X _08012_/Y _08010_/X _08009_/X _10059_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_13508__625 VPWR VGND VPWR VGND _14783_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
Xhold611 hold611/X hold611/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold600 hold600/X hold600/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 hold622/X hold622/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 hold633/X hold633/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 hold644/X hold644/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 hold666/X hold666/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold677 hold677/X hold677/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 hold655/X hold655/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold688/X hold688/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 hold699/X hold699/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ VPWR VGND VGND VPWR _12846_/B _12845_/B _15571_/Q sky130_fd_sc_hd__nor2_2
X_09895_ VPWR VGND VPWR VGND _15480_/Q hold1442/X _09907_/S _09895_/X sky130_fd_sc_hd__a21o_1
X_08915_ VGND VPWR VGND VPWR _15135_/D hold1241/X _08919_/A2 _08914_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
Xhold1300 hold1300/X _14848_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 hold1322/X _14128_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14112__1229 VPWR VGND VPWR VGND _15531_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
Xhold1333 hold1333/X _15626_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1311 _15607_/D _09981_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ VGND VPWR VPWR VGND _15167_/D _09689_/A0 _08846_/S hold609/X sky130_fd_sc_hd__mux2_1
Xhold1344 hold1344/X _15347_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1366 _10028_/A _15627_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1355 _10035_/A _15630_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 hold1377/X _15068_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_849 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08777_ VGND VPWR VPWR VGND _15229_/D _09726_/A1 _08779_/S hold215/X sky130_fd_sc_hd__mux2_1
Xhold1388 _08379_/A _15397_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 _08818_/A _15194_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13060__177 VPWR VGND VPWR VGND _14303_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07728_ VPWR VGND VGND VPWR _07794_/B _15559_/Q _07728_/B sky130_fd_sc_hd__or2_1
X_07659_ VPWR VGND VPWR VGND _07659_/B _07659_/C _07659_/A _07659_/X sky130_fd_sc_hd__or3_4
XFILLER_41_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_43_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10670_ VGND VPWR VPWR VGND _10670_/X hold756/A _10670_/S hold166/A sky130_fd_sc_hd__mux2_1
X_09329_ VGND VPWR VPWR VGND _14715_/D hold409/X _09336_/S fanout33/X sky130_fd_sc_hd__mux2_1
Xclone44 VPWR VGND clone44/X clone44/A VPWR VGND sky130_fd_sc_hd__buf_6
X_12340_ VGND VPWR VGND VPWR _12340_/X _15019_/Q _12705_/A2 _12591_/S _12339_/X sky130_fd_sc_hd__o211a_1
Xclone55 VGND VPWR clone55/X clone55/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_12271_ VGND VPWR VPWR VGND _12275_/B _14622_/Q _12701_/S _14654_/Q sky130_fd_sc_hd__mux2_1
X_11222_ VGND VPWR VGND VPWR _11222_/X _11219_/X _11221_/X _10816_/A _11259_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_0_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11153_ VPWR VGND _11153_/X _11152_/X _11148_/X _11246_/S _11144_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11084_ VGND VPWR VPWR VGND _11084_/X _11083_/X _11092_/S _11082_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10104_ VPWR VGND VGND VPWR _10104_/X hold369/A _10609_/S sky130_fd_sc_hd__or2_1
X_14912_ hold581/A _14912_/CLK _14912_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10035_ VPWR VGND VGND VPWR _10035_/A _10035_/B _10036_/B sky130_fd_sc_hd__nor2_1
X_14843_ _14843_/Q clkload19/A _14843_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13301__418 VPWR VGND VPWR VGND _14576_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_14774_ hold605/A _14774_/CLK _14774_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11986_ VGND VPWR VPWR VGND _11986_/X hold631/A _11998_/S hold284/A sky130_fd_sc_hd__mux2_1
X_10937_ VGND VPWR VPWR VGND _10937_/X hold603/A _11179_/S hold336/A sky130_fd_sc_hd__mux2_1
XFILLER_32_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_16_286 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10868_ VGND VPWR VPWR VGND _10868_/X _14208_/Q _10885_/S _15216_/Q sky130_fd_sc_hd__mux2_1
X_12607_ VGND VPWR VPWR VGND _12607_/X hold456/A _12623_/S hold326/A sky130_fd_sc_hd__mux2_1
X_10799_ VGND VPWR VGND VPWR _10799_/X hold790/A _11215_/A2 _10798_/X _11213_/S sky130_fd_sc_hd__o211a_1
X_15326_ _15326_/Q _15326_/CLK _15326_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12538_ VGND VPWR VPWR VGND _12542_/B hold641/A _12539_/S hold283/A sky130_fd_sc_hd__mux2_1
XFILLER_8_452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15257_ hold553/A _15257_/CLK _15257_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12469_ VGND VPWR VGND VPWR _12469_/X _12489_/A1 _12465_/X _12468_/X _12485_/C1 sky130_fd_sc_hd__o211a_1
X_14208_ _14208_/Q _14208_/CLK _14208_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15188_ hold775/A _15188_/CLK _15188_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14139_ _14139_/Q _14139_/CLK _14139_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout409 VPWR VGND _10622_/C1 _08178_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
X_08700_ VGND VPWR VGND VPWR _08700_/X _08700_/A2 _08700_/B1 _15280_/Q _08699_/X sky130_fd_sc_hd__a211o_1
X_09680_ VGND VPWR VPWR VGND _14360_/D hold857/X _09684_/S fanout21/X sky130_fd_sc_hd__mux2_1
X_08631_ VPWR VGND VGND VPWR _08630_/X _08690_/S _08194_/Y _14410_/Q _08631_/X _08629_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_687 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_55_849 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_54_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08562_ VPWR VGND VGND VPWR _08562_/A _08980_/B _08562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_78_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08493_ VPWR VGND VGND VPWR _08522_/B _14766_/Q _08493_/Y sky130_fd_sc_hd__nand2b_1
X_07513_ VPWR VGND VPWR VGND _07547_/B _07547_/A _07547_/C _07513_/X sky130_fd_sc_hd__a21o_1
X_07444_ VPWR VGND VPWR VGND _08548_/A _08559_/A _08554_/A _08566_/A _07444_/X sky130_fd_sc_hd__or4_1
Xfanout38 VGND VPWR _07953_/X fanout38/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout16 VGND VPWR _08070_/X fanout16/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_35_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout27 VGND VPWR fanout28/X fanout27/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_22_212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout49 VPWR VGND fanout49/X _07890_/X VPWR VGND sky130_fd_sc_hd__buf_6
X_07375_ VGND VPWR VGND VPWR _08081_/A _08137_/C _08137_/A _08137_/B _08116_/A sky130_fd_sc_hd__a211o_1
X_13916__1033 VPWR VGND VPWR VGND _15288_/CLK clkload50/A sky130_fd_sc_hd__inv_2
X_09114_ VGND VPWR VPWR VGND _14981_/D hold331/X _09128_/S fanout25/X sky130_fd_sc_hd__mux2_1
X_09045_ VGND VPWR VPWR VGND _15045_/D hold736/X _09059_/S fanout25/X sky130_fd_sc_hd__mux2_1
XFILLER_11_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13742__859 VPWR VGND VPWR VGND _15114_/CLK clkload46/A sky130_fd_sc_hd__inv_2
Xhold452 hold452/X hold452/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 hold463/X hold463/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 hold430/X hold430/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 hold441/X hold441/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12971__88 VPWR VGND VPWR VGND _14214_/CLK clkload52/A sky130_fd_sc_hd__inv_2
Xhold485 hold485/X hold485/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 hold474/X hold474/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold496/X hold496/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09947_ VPWR VGND VPWR VGND _14128_/Q _09947_/C _14129_/Q _09954_/C sky130_fd_sc_hd__or3_1
X_13595__712 VPWR VGND VPWR VGND _14935_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_09878_ VPWR VGND VGND VPWR _09878_/A _09878_/Y _09878_/B sky130_fd_sc_hd__nand2_1
Xhold1130 _11555_/A _15438_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 hold1141/X _15250_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 _11561_/A _15441_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1152 hold1152/X _14139_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ VGND VPWR VPWR VGND _08847_/S fanout48/X hold1219/X _15184_/D sky130_fd_sc_hd__mux2_2
Xhold1185 hold1185/X _14686_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 hold1163/X _14174_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13636__753 VPWR VGND VPWR VGND _14976_/CLK clkload13/A sky130_fd_sc_hd__inv_2
Xhold1196 hold1196/X _15502_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_808 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11840_ VGND VPWR VGND VPWR _11840_/X _11958_/A _11836_/X _11839_/X _12184_/C1 sky130_fd_sc_hd__o211a_1
X_11771_ VGND VPWR VPWR VGND _11771_/X hold816/A _12006_/B hold671/A sky130_fd_sc_hd__mux2_1
X_10722_ VGND VPWR VPWR VGND _10722_/X _14204_/Q _10743_/B hold550/A sky130_fd_sc_hd__mux2_1
X_14490_ hold996/A _14490_/CLK _14490_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_216 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10653_ VPWR VGND VPWR VGND _10652_/X _10667_/C1 _10651_/X _10653_/Y sky130_fd_sc_hd__a21oi_1
X_10584_ VGND VPWR VPWR VGND _10584_/X hold894/A _10730_/S hold298/A sky130_fd_sc_hd__mux2_1
X_15111_ _15111_/Q _15111_/CLK _15111_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12323_ VPWR VGND VPWR VGND _12322_/X _12703_/A1 _12321_/X _12323_/Y sky130_fd_sc_hd__a21oi_1
Xclkload19 clkload19/Y clkload19/A VGND VPWR VGND VPWR sky130_fd_sc_hd__clkinv_16
X_15042_ hold796/A _15042_/CLK _15042_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12254_ VPWR VGND VGND VPWR _12254_/X _12256_/S _12254_/B sky130_fd_sc_hd__or2_1
XFILLER_79_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11205_ VPWR VGND VGND VPWR _11205_/X _11205_/A _11205_/B sky130_fd_sc_hd__or2_1
X_12185_ VGND VPWR VGND VPWR _12185_/X _12185_/A1 _12180_/X _12184_/X _12222_/C1 sky130_fd_sc_hd__o211a_1
X_11136_ VPWR VGND VGND VPWR _11173_/A _11136_/B _11136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_694 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11067_ VGND VPWR VGND VPWR _11067_/X hold738/A _11184_/A2 _11066_/X _11178_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10018_ VPWR VGND VPWR VGND _10017_/C _15622_/Q hold1278/X _10019_/B sky130_fd_sc_hd__a21oi_1
X_14826_ _14826_/Q clkload30/A _14826_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13379__496 VPWR VGND VPWR VGND _14654_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
XFILLER_52_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_75_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14757_ hold296/A _14757_/CLK _14757_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11969_ VPWR VGND VPWR VGND _11968_/X _11966_/X _11967_/X _11969_/X _12175_/A1 sky130_fd_sc_hd__a22o_1
XFILLER_36_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14688_ hold697/A _14688_/CLK _14688_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14203__921 _14203_/D _14203__921/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_07160_ VPWR VGND VGND VPWR _14407_/Q _07301_/A2 _07301_/B1 _07162_/B sky130_fd_sc_hd__o21a_1
X_14111__1228 VPWR VGND VPWR VGND _15530_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_15309_ hold989/A _15309_/CLK _15309_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07091_ VPWR VGND VPWR VGND _11899_/A _15453_/Q sky130_fd_sc_hd__inv_2
XFILLER_8_271 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout217 VPWR VGND fanout217/X _07978_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout206 VGND VPWR _12375_/S _12489_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout228 VGND VPWR _12739_/C1 _12662_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09801_ VPWR VGND VGND VPWR _09801_/X _09801_/A _09827_/S sky130_fd_sc_hd__or2_1
Xfanout239 VGND VPWR _08270_/A1 _12193_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13323__440 VPWR VGND VPWR VGND _14598_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07993_ VPWR VGND VGND VPWR _07993_/A _07993_/B _07994_/C sky130_fd_sc_hd__nor2_1
X_09732_ _14314_/D fanout91/X fanout87/X _09730_/Y _09731_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xtt_um_femto_900 uio_out[3] tt_um_femto_900/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09663_ VGND VPWR VPWR VGND _14377_/D hold980/X _09675_/S fanout86/X sky130_fd_sc_hd__mux2_1
X_08614_ VPWR VGND VGND VPWR _08617_/A _09007_/B _08614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09594_ _14474_/D fanout92/X fanout88/X _09592_/Y _09593_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08545_ VPWR VGND VGND VPWR _08545_/A _08546_/B _08559_/B sky130_fd_sc_hd__nand2_1
X_08476_ VPWR VGND VGND VPWR _08476_/X _08476_/A _08482_/B sky130_fd_sc_hd__or2_1
X_07427_ VPWR VGND VGND VPWR _15467_/Q _07429_/A _07519_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_1210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07358_ VPWR VGND VGND VPWR _11899_/A _07358_/B _08117_/B sky130_fd_sc_hd__nor2_1
X_13172__289 VPWR VGND VPWR VGND _14447_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_10_237 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_40_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07289_ VGND VPWR VGND VPWR _07286_/B _07926_/A _07946_/A _07811_/B sky130_fd_sc_hd__o21ba_1
X_09028_ _15062_/D fanout93/X fanout89/X _09055_/S _09027_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_46_1003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold271 hold271/X hold271/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold260 hold260/X hold260/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/X hold282/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/X hold293/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout751 VPWR VGND _12822_/A _12789_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout740 VPWR VGND _11537_/S _09965_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout762 VPWR VGND _08249_/A2 _08002_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout773 VGND VPWR _08066_/B _07859_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout784 VGND VPWR _07304_/A2 _07301_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13066__183 VPWR VGND VPWR VGND _14309_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
XFILLER_74_911 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout795 VGND VPWR _08700_/A2 _08667_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_12872_ VGND VPWR VPWR VGND _15596_/D _07661_/X _14802_/D _15596_/Q sky130_fd_sc_hd__mux2_1
XFILLER_46_668 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_100 _12740_/C1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_34_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13870__987 VPWR VGND VPWR VGND _15242_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_14611_ hold806/A _14611_/CLK _14611_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11823_ VGND VPWR VGND VPWR _11823_/X _11820_/X _11822_/X _12748_/A1 _12744_/C1 sky130_fd_sc_hd__a211o_1
XANTENNA_122 _10893_/B1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_111 clone2/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_57_1121 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15591_ _15591_/Q clkload49/A _15591_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14542_ hold503/A _14542_/CLK _14542_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11754_ VGND VPWR VPWR VGND _11754_/X hold864/A _12094_/S hold395/A sky130_fd_sc_hd__mux2_1
X_14473_ hold604/A _14473_/CLK _14473_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10705_ VPWR VGND VGND VPWR _10705_/X _10705_/A _10705_/B sky130_fd_sc_hd__or2_1
XFILLER_35_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11685_ VGND VPWR VPWR VGND _11685_/X _11682_/X _12476_/S _11681_/X sky130_fd_sc_hd__mux2_1
X_10636_ VPWR VGND VPWR VGND _10635_/X _10618_/A _12121_/B1 _10636_/X sky130_fd_sc_hd__a21o_1
X_13764__881 VPWR VGND VPWR VGND _15136_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_10567_ VGND VPWR VPWR VGND _10567_/X hold640/A _10567_/S hold260/A sky130_fd_sc_hd__mux2_1
XFILLER_6_742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12306_ VPWR VGND VPWR VGND _12305_/X _12584_/A _12602_/B1 _12306_/X sky130_fd_sc_hd__a21o_1
X_10498_ VGND VPWR VPWR VGND _10502_/B hold601/A _10516_/S hold360/A sky130_fd_sc_hd__mux2_1
X_12237_ VGND VPWR VGND VPWR _12237_/X _12234_/X _12236_/X _12256_/S _12596_/C1 sky130_fd_sc_hd__a211o_1
X_15025_ _15025_/Q _15025_/CLK _15025_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13307__424 VPWR VGND VPWR VGND _14582_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_12168_ VGND VPWR VPWR VGND _12172_/B hold608/A _12171_/S hold185/A sky130_fd_sc_hd__mux2_1
XFILLER_2_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11119_ VGND VPWR VPWR VGND _11123_/B hold629/A _11142_/S hold388/A sky130_fd_sc_hd__mux2_1
X_12099_ VGND VPWR VGND VPWR _12099_/X _12099_/A1 _12095_/X _12098_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
X_13915__1032 VPWR VGND VPWR VGND _15287_/CLK clkload50/A sky130_fd_sc_hd__inv_2
XFILLER_37_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14809_ hold153/A _14809_/CLK _14809_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_45_690 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08330_ VGND VPWR VPWR VGND _15489_/D _09547_/A1 _08330_/S hold821/X sky130_fd_sc_hd__mux2_1
X_08261_ VPWR VGND VGND VPWR _15447_/Q _07222_/A _08278_/B _08261_/X sky130_fd_sc_hd__o21a_1
X_07212_ VGND VPWR VPWR VGND _07220_/S _15595_/Q _14384_/Q _07369_/B sky130_fd_sc_hd__mux2_2
X_08192_ VPWR VGND VPWR VGND _08174_/Y _15337_/Q _08491_/A _08192_/X _14840_/Q sky130_fd_sc_hd__a22o_1
X_07143_ VPWR VGND VPWR VGND wire858/A _07143_/A1 _08294_/B1 _07143_/X _12878_/A sky130_fd_sc_hd__a22o_1
X_12941__58 VPWR VGND VPWR VGND _14184_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_07976_ VPWR VGND VPWR VGND _07976_/X _07976_/A _07976_/B sky130_fd_sc_hd__or2_2
XFILLER_28_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09715_ VGND VPWR VPWR VGND _14328_/D fanout20/X _09721_/S hold752/X sky130_fd_sc_hd__mux2_1
X_09646_ VGND VPWR VPWR VGND _14424_/D hold898/X _09657_/S fanout20/X sky130_fd_sc_hd__mux2_1
XFILLER_56_977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_35_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13100__217 VPWR VGND VPWR VGND _14343_/CLK clkload42/A sky130_fd_sc_hd__inv_2
XFILLER_58_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09577_ VGND VPWR VPWR VGND _14488_/D hold906/X _09588_/S fanout19/X sky130_fd_sc_hd__mux2_1
X_08528_ VPWR VGND VPWR VGND _08540_/B1 hold1444/X _08503_/A _08529_/B _15322_/Q sky130_fd_sc_hd__a22o_1
XFILLER_19_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08459_ VGND VPWR VGND VPWR _15347_/D hold1108/X _08458_/B _08458_/Y _08919_/C1 sky130_fd_sc_hd__o211a_1
X_13748__865 VPWR VGND VPWR VGND _15120_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_1062 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11470_ VGND VPWR VPWR VGND _11470_/X _11469_/X _11476_/S _15454_/Q sky130_fd_sc_hd__mux2_1
X_10421_ VGND VPWR VPWR VGND _10421_/X hold455/A _10720_/S hold330/A sky130_fd_sc_hd__mux2_1
X_10352_ VGND VPWR VPWR VGND _10352_/X _14194_/Q _10353_/S hold225/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12022_ VGND VPWR VPWR VGND _12022_/X _14199_/Q _12190_/S hold324/A sky130_fd_sc_hd__mux2_1
X_10283_ VPWR VGND VPWR VGND _10282_/X _10608_/A1 _10281_/X _10283_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout581 VPWR VGND _09272_/S _09241_/Y VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout570 _09414_/S _09406_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_19_624 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout592 VGND VPWR _08816_/Y _08842_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_14110__1227 VPWR VGND VPWR VGND _15529_/CLK clkload20/A sky130_fd_sc_hd__inv_2
XFILLER_73_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12855_ VGND VPWR VPWR VGND _15579_/D _08112_/Y _12877_/S _12855_/A0 sky130_fd_sc_hd__mux2_1
X_11806_ VGND VPWR VPWR VGND _11807_/B _11805_/Y _12583_/S _11797_/Y sky130_fd_sc_hd__mux2_1
X_15574_ _15574_/Q clkload32/A _15574_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12786_ VPWR VGND VGND VPWR _10079_/X _08078_/Y _12788_/S _08076_/Y _12786_/X _12785_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14525_ hold311/A _14525_/CLK _14525_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11737_ VPWR VGND VGND VPWR _11737_/X hold578/A _12409_/B sky130_fd_sc_hd__or2_1
X_11668_ VGND VPWR VPWR VGND _11668_/X hold426/A _11965_/S hold355/A sky130_fd_sc_hd__mux2_1
X_14456_ hold744/A _14456_/CLK _14456_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14387_ _14387_/Q clkload21/A _14387_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11599_ VPWR VGND VGND VPWR _11599_/X hold192/A _11998_/S sky130_fd_sc_hd__or2_1
X_10619_ VPWR VGND VGND VPWR _10619_/X hold488/A _10627_/S sky130_fd_sc_hd__or2_1
XFILLER_6_550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15008_ _15008_/Q _15008_/CLK _15008_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13541__658 VPWR VGND VPWR VGND _14872_/CLK clkload24/A sky130_fd_sc_hd__inv_2
XFILLER_57_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07830_ VGND VPWR _08220_/B _15546_/Q _15547_/Q _15545_/Q VPWR VGND sky130_fd_sc_hd__and3_1
X_07761_ VPWR VGND VGND VPWR _07759_/X _07761_/B _08218_/A sky130_fd_sc_hd__nand2b_1
X_13394__511 VPWR VGND VPWR VGND _14669_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_09500_ VGND VPWR VPWR VGND _14559_/D fanout47/X _09514_/S hold571/X sky130_fd_sc_hd__mux2_1
XFILLER_65_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07692_ VPWR VGND VPWR VGND _10893_/B1 _07119_/A clone17/A _07692_/Y sky130_fd_sc_hd__a21oi_1
X_09431_ VGND VPWR VPWR VGND _14621_/D fanout39/X _09443_/S hold619/X sky130_fd_sc_hd__mux2_1
XFILLER_53_936 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09362_ VGND VPWR VPWR VGND _14684_/D hold722/X _09377_/S fanout36/X sky130_fd_sc_hd__mux2_1
X_13435__552 VPWR VGND VPWR VGND _14710_/CLK clkload11/A sky130_fd_sc_hd__inv_2
X_08313_ VGND VPWR VPWR VGND _15506_/D fanout64/X _08318_/S hold914/X sky130_fd_sc_hd__mux2_1
XANTENNA_22 _14389_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_09293_ VGND VPWR VPWR VGND _14748_/D fanout35/X _09302_/S hold211/X sky130_fd_sc_hd__mux2_1
XANTENNA_11 _08212_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_44 fanout282/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_66 _08806_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_55 _12080_/A2 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08244_ VPWR VGND VPWR VGND _15068_/Q _08293_/B1 _08244_/X _08263_/A2 _07219_/X _08243_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_33 _12373_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_99 fanout234/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08175_ VPWR VGND VPWR VGND _08174_/Y _15338_/Q _08491_/A _08175_/X _14841_/Q sky130_fd_sc_hd__a22o_1
XANTENNA_88 _14383_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_77 _08366_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07126_ VPWR VGND VPWR VGND _07126_/Y _14842_/Q sky130_fd_sc_hd__inv_2
X_07959_ _07959_/X _07800_/B _07959_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_10970_ VPWR VGND VGND VPWR _10951_/Y _10969_/X _12677_/A2 _14402_/Q _14402_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_09629_ VGND VPWR VPWR VGND _14441_/D hold934/X _09637_/S fanout86/X sky130_fd_sc_hd__mux2_1
X_12640_ VPWR VGND VGND VPWR _12621_/Y _12639_/X _12677_/A2 _15473_/Q _15473_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_13178__295 VPWR VGND VPWR VGND _14453_/CLK clkload24/A sky130_fd_sc_hd__inv_2
XFILLER_58_1282 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_1233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12571_ VPWR VGND VGND VPWR _12571_/X _12581_/S _12571_/B sky130_fd_sc_hd__or2_1
X_14310_ _14310_/Q _14310_/CLK _14310_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_50_clk clkload42/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_11_332 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11522_ VGND VPWR VPWR VGND _15091_/D _11521_/X _11528_/S _15091_/Q sky130_fd_sc_hd__mux2_1
X_15290_ _15290_/Q _15290_/CLK _15290_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_354 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11453_ VGND VPWR VPWR VGND _15068_/D _11452_/X _11480_/S hold1377/X sky130_fd_sc_hd__mux2_1
X_14241_ _14241_/Q _14241_/CLK _14241_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10404_ VGND VPWR VGND VPWR _10404_/X _10693_/B1 _10399_/X _10403_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_13914__1031 VPWR VGND VPWR VGND _15286_/CLK clkload50/A sky130_fd_sc_hd__inv_2
X_14172_ hold422/A _14172_/CLK _14172_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11384_ VGND VPWR VPWR VGND _11384_/X _11383_/X _11387_/S _14849_/Q sky130_fd_sc_hd__mux2_1
X_10335_ VPWR VGND VGND VPWR _10335_/X _11112_/A _10335_/B sky130_fd_sc_hd__or2_1
XFILLER_3_531 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10266_ VPWR VGND VPWR VGND _10265_/X _11210_/A _12491_/B1 _10266_/X sky130_fd_sc_hd__a21o_1
X_12005_ VGND VPWR VPWR VGND _12005_/X hold367/A _12005_/S hold796/A sky130_fd_sc_hd__mux2_1
X_13876__993 VPWR VGND VPWR VGND _15248_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_10197_ VGND VPWR VPWR VGND _10197_/X hold503/A _10567_/S hold219/A sky130_fd_sc_hd__mux2_1
Xclone146 VPWR VGND clone146/X fanout79/X VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_19_410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13419__536 VPWR VGND VPWR VGND _14694_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_15626_ _15626_/Q clkload49/A _15626_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12838_ VPWR VGND VGND VPWR _12837_/X _09961_/Y _11458_/S _07360_/B _15568_/D _11477_/S
+ sky130_fd_sc_hd__o221a_1
X_12769_ VPWR VGND VPWR VGND _08157_/B _12817_/A _12878_/C _12769_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_41_clk clkload49/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_15557_ _15557_/Q clkload43/A _15557_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15488_ _15488_/Q _15488_/CLK _15488_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14508_ hold250/A _14508_/CLK _14508_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14439_ hold941/A _14439_/CLK _14439_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold837 hold837/X hold837/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 hold826/X hold826/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold804 hold804/X hold804/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 hold815/X hold815/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ VPWR VGND VPWR VGND _09979_/X _09909_/A _09938_/A _14767_/D sky130_fd_sc_hd__a21oi_1
X_12986__103 VPWR VGND VPWR VGND _14229_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
Xhold859 hold859/X hold859/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 hold848/X hold848/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08931_ VGND VPWR _09892_/A _15162_/Q _09890_/A _09970_/B VPWR VGND sky130_fd_sc_hd__and3_1
X_12911__28 VPWR VGND VPWR VGND _14154_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_08862_ VGND VPWR _08868_/B _15480_/Q _15162_/Q _08862_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_07813_ VPWR VGND VGND VPWR _07813_/A _07813_/B _07854_/B sky130_fd_sc_hd__nor2_1
X_08793_ VGND VPWR VPWR VGND _08811_/S fanout48/X hold1131/X _15216_/D sky130_fd_sc_hd__mux2_2
X_07744_ VPWR VGND VPWR VGND _07751_/C _11535_/A _15553_/Q _08096_/A sky130_fd_sc_hd__a21oi_1
X_07675_ VGND VPWR VGND VPWR _15357_/Q _07558_/B _15130_/Q _07676_/A clone18/X sky130_fd_sc_hd__a22oi_4
XFILLER_16_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_77_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09414_ VGND VPWR VPWR VGND _14635_/D hold692/X _09414_/S fanout97/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clkload48/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09345_ VGND VPWR VPWR VGND _14699_/D hold531/X _09345_/S fanout95/X sky130_fd_sc_hd__mux2_1
X_09276_ VPWR VGND VGND VPWR _09729_/A _09276_/Y _09591_/A sky130_fd_sc_hd__nor2_2
X_08227_ VPWR VGND VPWR VGND _15069_/Q _08293_/B1 _08227_/X _08263_/A2 _07216_/X _08226_/X
+ sky130_fd_sc_hd__a221o_1
X_13212__329 VPWR VGND VPWR VGND _14487_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_08158_ VPWR VGND VGND VPWR _08201_/C _08223_/A _08223_/B sky130_fd_sc_hd__or2_1
X_07109_ VPWR VGND VPWR VGND _07109_/Y _14819_/Q sky130_fd_sc_hd__inv_2
X_08089_ VPWR VGND VGND VPWR _08220_/A _08076_/Y _08147_/A _08078_/Y _08089_/X sky130_fd_sc_hd__o22a_1
X_13563__680 VPWR VGND VPWR VGND _14894_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_10120_ VGND VPWR VPWR VGND _10124_/B hold519/A _10612_/S hold460/A sky130_fd_sc_hd__mux2_1
X_10051_ VGND VPWR _10051_/B _10051_/Y _10051_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13106__223 VPWR VGND VPWR VGND _14349_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
XFILLER_25_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14790_ _14790_/Q _14790_/CLK _14790_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10953_ VGND VPWR VPWR VGND _10953_/X hold866/A _11179_/S hold454/A sky130_fd_sc_hd__mux2_1
X_10884_ VGND VPWR VPWR VGND _10888_/B _15184_/Q _10885_/S hold707/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_clk clkload30/A clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_31_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12623_ VGND VPWR VPWR VGND _12623_/X hold793/A _12623_/S hold598/A sky130_fd_sc_hd__mux2_1
X_15411_ hold437/A _15411_/CLK _15411_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15342_ _15342_/Q _15342_/CLK _15342_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12554_ VGND VPWR VPWR VGND _12554_/X _12553_/X _12665_/S _12552_/X sky130_fd_sc_hd__mux2_1
X_11505_ VGND VPWR VPWR VGND _11505_/X _15087_/Q _11535_/C _15085_/Q sky130_fd_sc_hd__mux2_1
X_15273_ hold840/A _15273_/CLK _15273_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12977__94 VPWR VGND VPWR VGND _14220_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_14224_ hold229/A _14224_/CLK _14224_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12485_ VGND VPWR VGND VPWR _12485_/X _12482_/X _12484_/X _12489_/A1 _12485_/C1 sky130_fd_sc_hd__a211o_1
X_11436_ VGND VPWR VGND VPWR _11436_/X _14933_/Q _07109_/Y _11439_/A2 sky130_fd_sc_hd__a21bo_1
X_13804__921 VPWR VGND VPWR VGND _15176_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_11367_ VGND VPWR _14854_/Q _14852_/Q _11368_/C _11367_/D _14851_/Q VPWR VGND sky130_fd_sc_hd__and4b_1
XFILLER_4_851 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14155_ hold625/A _14155_/CLK _14155_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10318_ VGND VPWR VGND VPWR _10318_/X _14257_/Q _11262_/A2 _10317_/X _10315_/S sky130_fd_sc_hd__o211a_1
X_11298_ VPWR VGND _14817_/D _11298_/B _11388_/S VPWR VGND sky130_fd_sc_hd__and2_1
X_10249_ VPWR VGND VGND VPWR _10249_/X hold556/A _10924_/B sky130_fd_sc_hd__or2_1
XFILLER_78_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14988_ hold748/A _14988_/CLK _14988_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_755 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_23_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07460_ VPWR VGND VGND VPWR _15451_/Q _07462_/A _15596_/Q sky130_fd_sc_hd__nand2_1
X_15609_ _15609_/Q clkload27/A _15609_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07391_ _07391_/X _07292_/B _15468_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_14_clk clkload22/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09130_ VPWR VGND VPWR VGND _09130_/Y _09157_/S sky130_fd_sc_hd__inv_2
X_09061_ VPWR VGND VPWR VGND _09061_/X _09095_/B _09764_/A sky130_fd_sc_hd__or2_2
X_08012_ VPWR VGND VPWR VGND _10072_/B _15080_/Q _08011_/X _08012_/Y sky130_fd_sc_hd__a21oi_1
X_13547__664 VPWR VGND VPWR VGND _14878_/CLK clkload21/A sky130_fd_sc_hd__inv_2
Xhold601 hold601/X hold601/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 hold612/X hold612/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 hold645/X hold645/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 hold623/X hold623/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 hold634/X hold634/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ VPWR VGND VGND VPWR _12846_/B _15570_/Q _12842_/B sky130_fd_sc_hd__or2_1
Xhold678 hold678/X hold678/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold667 hold667/X hold667/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 hold656/X hold656/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ VPWR VGND VGND VPWR _08914_/X _08914_/A _08926_/B sky130_fd_sc_hd__or2_1
Xhold689 hold689/X hold689/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09894_ VGND VPWR VPWR VGND _14146_/D _09907_/S _09894_/S _09893_/Y sky130_fd_sc_hd__mux2_1
Xhold1312 hold1312/X _14844_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1334 _10026_/B _10025_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 _09995_/A _15613_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1301 hold1301/X _15620_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ VGND VPWR VPWR VGND _15168_/D _09550_/A1 _08850_/S hold523/X sky130_fd_sc_hd__mux2_1
Xhold1345 hold1345/X _14934_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1367 hold1367/X _15360_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08776_ VGND VPWR VPWR VGND _15230_/D _09864_/A0 _08776_/S hold484/X sky130_fd_sc_hd__mux2_1
XFILLER_22_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1356 _08747_/A _15258_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07727_ VPWR VGND _07727_/X _07728_/B _15559_/Q VPWR VGND sky130_fd_sc_hd__and2_1
Xhold1378 hold1378/X _14378_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13913__1030 VPWR VGND VPWR VGND _15285_/CLK clkload16/A sky130_fd_sc_hd__inv_2
XFILLER_27_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1389 _09696_/A _14346_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07658_ _07659_/C _07655_/X _07656_/X _07657_/X _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07589_ VGND VPWR VGND VPWR _08491_/A _08174_/A _07588_/X _07589_/X _15339_/Q sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09328_ VGND VPWR VPWR VGND _14716_/D hold418/X _09336_/S fanout36/X sky130_fd_sc_hd__mux2_1
X_09259_ VGND VPWR VPWR VGND _14784_/D fanout31/X _09275_/S hold608/X sky130_fd_sc_hd__mux2_1
Xclone45 VGND VPWR clone45/X clone45/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_12270_ VGND VPWR VGND VPWR _15463_/D _12602_/B1 _12268_/X _12269_/X _11341_/A sky130_fd_sc_hd__o211a_1
X_11221_ VGND VPWR VGND VPWR _11221_/X hold814/A _11262_/A2 _11220_/X _10851_/A sky130_fd_sc_hd__o211a_1
XFILLER_4_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11152_ VGND VPWR VGND VPWR _11152_/X _11149_/X _11151_/X _11189_/A1 _11245_/A1 sky130_fd_sc_hd__a211o_1
X_10103_ VGND VPWR VPWR VGND _10103_/X _10102_/X _10144_/S _10101_/X sky130_fd_sc_hd__mux2_1
X_11083_ VGND VPWR VPWR VGND _11083_/X _14502_/Q _11091_/S _14182_/Q sky130_fd_sc_hd__mux2_1
XFILLER_66_1381 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_803 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10034_ VPWR VGND _10038_/C _10035_/B _15630_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_7_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14911_ hold466/A _14911_/CLK _14911_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14842_ _14842_/Q clkload30/A _14842_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13340__457 VPWR VGND VPWR VGND _14615_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_14773_ hold534/A _14773_/CLK _14773_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11985_ VGND VPWR VPWR VGND _11985_/X _14198_/Q _11998_/S hold341/A sky130_fd_sc_hd__mux2_1
X_10936_ VGND VPWR VPWR VGND _10936_/X hold713/A _11179_/S _15250_/Q sky130_fd_sc_hd__mux2_1
X_13193__310 VPWR VGND VPWR VGND _14468_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_10867_ VGND VPWR VGND VPWR _10867_/X _10891_/C1 _10862_/X _10866_/X _12869_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_44_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12606_ VGND VPWR VPWR VGND _12606_/X hold564/A _12623_/S hold348/A sky130_fd_sc_hd__mux2_1
X_13234__351 VPWR VGND VPWR VGND _14509_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_10798_ VPWR VGND VGND VPWR _10798_/X _14302_/Q _11204_/S sky130_fd_sc_hd__or2_1
X_15325_ hold923/A _15325_/CLK hold924/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12537_ VPWR VGND VPWR VGND _12536_/X _12656_/A1 _12535_/X _12537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_987 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12468_ VPWR VGND VGND VPWR _12468_/X _12470_/S _12468_/B sky130_fd_sc_hd__or2_1
X_15256_ hold247/A _15256_/CLK _15256_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11419_ VPWR VGND VPWR VGND _11418_/X _11417_/X _09938_/A _14860_/D sky130_fd_sc_hd__a21o_1
X_14207_ _14207_/Q _14207_/CLK _14207_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15187_ hold416/A _15187_/CLK _15187_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14138_ _14138_/Q _14138_/CLK _14138_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12399_ VPWR VGND VGND VPWR _12732_/A _12399_/B _12399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk clkload8/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_80_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08630_ VPWR VGND VGND VPWR _08630_/X _14394_/Q _08640_/B sky130_fd_sc_hd__or2_1
XFILLER_55_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08561_ VPWR VGND VPWR VGND _07736_/A _07523_/B _08980_/B _08559_/Y _08560_/X _07534_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_78_1285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08492_ _08492_/X _08522_/B _14766_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_07512_ VPWR VGND VGND VPWR _07512_/A _07547_/C _07512_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07443_ VPWR VGND VGND VPWR _08546_/A _08559_/A _08545_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout17 VPWR VGND fanout17/X _08070_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout28 VGND VPWR _08014_/X fanout28/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout39 VGND VPWR fanout40/X fanout39/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07374_ VPWR VGND VPWR VGND _08137_/C _08137_/B _08137_/A _08138_/A sky130_fd_sc_hd__a21oi_1
X_09113_ VGND VPWR VPWR VGND _14982_/D hold457/X _09126_/S fanout28/X sky130_fd_sc_hd__mux2_1
X_09044_ VGND VPWR VPWR VGND _15046_/D hold660/X _09051_/S _08014_/X sky130_fd_sc_hd__mux2_1
X_13781__898 VPWR VGND VPWR VGND _15153_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
Xhold420 hold420/X hold420/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 hold442/X hold442/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold431/X hold431/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 hold453/X hold453/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 hold475/X hold475/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 hold486/X hold486/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 hold464/X hold464/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ VPWR VGND VPWR VGND _09945_/Y hold1393/X _09956_/S _14129_/D _09937_/Y sky130_fd_sc_hd__a22o_1
Xhold497 hold497/X hold497/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_611 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09877_ VPWR VGND VGND VPWR _09877_/X _14150_/Q _09878_/B sky130_fd_sc_hd__or2_1
Xhold1131 hold1131/X _15216_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _09024_/B _15063_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1120 hold1120/X _14598_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1175 hold1175/X _14839_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 hold1164/X _15222_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13675__792 VPWR VGND VPWR VGND _15015_/CLK clkload20/A sky130_fd_sc_hd__inv_2
Xhold1153 hold1153/X _14184_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ VGND VPWR VPWR VGND _15185_/D fanout54/X _08846_/S hold428/X sky130_fd_sc_hd__mux2_1
X_08759_ VGND VPWR VPWR VGND _15247_/D fanout46/X _08773_/S hold317/X sky130_fd_sc_hd__mux2_1
Xhold1197 hold1197/X _15540_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 hold1186/X _15132_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11770_ VPWR VGND VGND VPWR _12103_/A _11770_/B _11770_/Y sky130_fd_sc_hd__nor2_1
X_10721_ VGND VPWR VPWR VGND _10721_/X hold544/A _10743_/B hold408/A sky130_fd_sc_hd__mux2_1
X_13218__335 VPWR VGND VPWR VGND _14493_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
XFILLER_70_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_41_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10652_ VGND VPWR VPWR VGND _10652_/X _10649_/X _10652_/S _10648_/X sky130_fd_sc_hd__mux2_1
X_10583_ VGND VPWR VGND VPWR _10583_/X _14875_/Q _10583_/A2 _10582_/X _10588_/S sky130_fd_sc_hd__o211a_1
X_15110_ hold954/A _15110_/CLK _15110_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12322_ VGND VPWR VPWR VGND _12322_/X _12319_/X _12684_/S _12318_/X sky130_fd_sc_hd__mux2_1
X_12947__64 VPWR VGND VPWR VGND _14190_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
XFILLER_68_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15041_ hold788/A _15041_/CLK _15041_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12253_ VGND VPWR VPWR VGND _12254_/B hold869/A _12578_/S hold742/A sky130_fd_sc_hd__mux2_1
XFILLER_5_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_68_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11204_ VGND VPWR VPWR VGND _11204_/X hold604/A _11204_/S hold249/A sky130_fd_sc_hd__mux2_1
X_12184_ VGND VPWR VGND VPWR _12184_/X _12183_/X _12182_/X _12164_/A _12184_/C1 sky130_fd_sc_hd__a211o_1
X_11135_ VGND VPWR VPWR VGND _11136_/B _11134_/Y _11246_/S _11126_/Y sky130_fd_sc_hd__mux2_1
XFILLER_49_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11066_ VPWR VGND VGND VPWR _11066_/X hold764/A _11175_/S sky130_fd_sc_hd__or2_1
XFILLER_1_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10017_ VGND VPWR _10021_/B _15623_/Q _15622_/Q _10017_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14825_ _14825_/Q clkload30/A _14825_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14756_ hold441/A _14756_/CLK _14756_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11968_ VGND VPWR VPWR VGND _11968_/X _11965_/X _11968_/S _11964_/X sky130_fd_sc_hd__mux2_1
X_14687_ hold565/A _14687_/CLK _14687_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11899_ VPWR VGND VGND VPWR _11899_/A _11899_/Y _11973_/B sky130_fd_sc_hd__nand2_1
X_10919_ VGND VPWR VPWR VGND _10919_/X hold987/A _10919_/S _14689_/Q sky130_fd_sc_hd__mux2_1
XFILLER_74_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15308_ hold865/A _15308_/CLK _15308_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07090_ VPWR VGND VPWR VGND _07376_/A _15454_/Q sky130_fd_sc_hd__inv_2
XFILLER_12_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15239_ hold187/A _15239_/CLK _15239_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13011__128 VPWR VGND VPWR VGND _14254_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_07992_ VGND VPWR _07992_/B _07993_/B _07992_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xfanout229 VGND VPWR _12739_/C1 _12670_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout218 VGND VPWR _12115_/C1 _12099_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout207 VGND VPWR _12375_/S _12720_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09800_ VPWR VGND VPWR VGND _09800_/Y _09827_/S sky130_fd_sc_hd__inv_2
X_09731_ VPWR VGND VGND VPWR _09731_/X _09731_/A _09757_/S sky130_fd_sc_hd__or2_1
X_13659__776 VPWR VGND VPWR VGND _14999_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Left_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xtt_um_femto_901 uio_out[4] tt_um_femto_901/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_39_154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09662_ _14378_/D fanout91/X fanout87/X _09687_/S _09661_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08613_ VGND VPWR VGND VPWR _15305_/D hold1063/X _08613_/A2 _08612_/X _09000_/C1
+ sky130_fd_sc_hd__o211a_1
X_09593_ VPWR VGND VGND VPWR _09593_/X _09593_/A _09622_/S sky130_fd_sc_hd__or2_1
XFILLER_78_1060 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08544_ VPWR VGND VGND VPWR _08559_/B _08544_/A _08544_/B sky130_fd_sc_hd__or2_1
XFILLER_78_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08475_ VGND VPWR VGND VPWR _15339_/D hold1233/X _08485_/A2 _08474_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_07426_ VGND VPWR VGND VPWR _07426_/X _07807_/S _07827_/C _15572_/Q _07703_/A sky130_fd_sc_hd__and4_2
XFILLER_39_1099 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07357_ VPWR VGND VPWR VGND _07356_/Y _07357_/Y _08083_/A _07196_/B sky130_fd_sc_hd__a21boi_1
XFILLER_17_1375 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09027_ VPWR VGND VGND VPWR hold1370/X _09055_/S _09027_/Y sky130_fd_sc_hd__nand2b_1
X_07288_ VPWR VGND VPWR VGND _07945_/A _07288_/A _07946_/A sky130_fd_sc_hd__or2_2
XFILLER_2_404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold261 hold261/X hold261/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13603__720 VPWR VGND VPWR VGND _14943_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_2_448 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold250 hold250/X hold250/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/X hold283/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/X hold272/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/X hold294/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout741 VGND VPWR _09965_/X _11530_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout730 VPWR VGND _10562_/B _11117_/B VPWR VGND sky130_fd_sc_hd__buf_4
X_09929_ VPWR VGND VPWR VGND _09928_/Y _14766_/Q _08522_/B _09929_/X _09912_/A sky130_fd_sc_hd__a22o_1
Xfanout763 VPWR VGND _07952_/A2 _07929_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout752 VPWR VGND _12789_/A _12831_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout785 VGND VPWR _07142_/X _07304_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout774 VPWR VGND _08066_/B _07415_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout796 VPWR VGND _08700_/A2 _08626_/A VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_4_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12871_ VGND VPWR VPWR VGND _15595_/D _07676_/Y _14802_/D _15595_/Q sky130_fd_sc_hd__mux2_1
XANTENNA_101 fanout314/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11822_ VGND VPWR VGND VPWR _11822_/X _15005_/Q _12746_/A2 _11810_/S _11821_/X sky130_fd_sc_hd__o211a_1
XANTENNA_112 _09825_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_14610_ hold462/A _14610_/CLK _14610_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_27_861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15590_ _15590_/Q clkload50/A _15590_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14541_ hold414/A _14541_/CLK _14541_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13452__569 VPWR VGND VPWR VGND _14727_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_11753_ VGND VPWR VPWR VGND _11757_/B hold784/A _12094_/S hold449/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10704_ VGND VPWR VGND VPWR _10704_/X _10705_/A _10700_/X _10703_/X _10704_/C1 sky130_fd_sc_hd__o211a_1
X_11684_ VGND VPWR VGND VPWR _11684_/X _12489_/A1 _11680_/X _11683_/X _12485_/C1 sky130_fd_sc_hd__o211a_1
X_14472_ hold656/A _14472_/CLK _14472_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10635_ VPWR VGND _10635_/X _10634_/X _10630_/X _10469_/S _10626_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12305_ VPWR VGND _12305_/X _12304_/X _12300_/X _12694_/S _12296_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_5_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10566_ VGND VPWR VPWR VGND _10566_/X hold752/A _10567_/S hold220/A sky130_fd_sc_hd__mux2_1
X_10497_ VPWR VGND VPWR VGND _10496_/X _10634_/C1 _10495_/X _10497_/Y sky130_fd_sc_hd__a21oi_1
X_12236_ VGND VPWR VGND VPWR _12236_/X _14493_/Q _12705_/A2 _12581_/S _12235_/X sky130_fd_sc_hd__o211a_1
X_15024_ _15024_/Q _15024_/CLK _15024_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13346__463 VPWR VGND VPWR VGND _14621_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_12167_ VPWR VGND VPWR VGND _12166_/X _12175_/A1 _12165_/X _12167_/Y sky130_fd_sc_hd__a21oi_1
X_11118_ VGND VPWR VGND VPWR _14406_/D _12602_/B1 _11116_/X _11117_/X _12751_/C1 sky130_fd_sc_hd__o211a_1
X_12098_ VPWR VGND VGND VPWR _12098_/X _12098_/A _12098_/B sky130_fd_sc_hd__or2_1
XFILLER_77_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11049_ VPWR VGND VGND VPWR _11049_/X _11176_/S _11049_/B sky130_fd_sc_hd__or2_1
X_14808_ _14808_/Q _14808_/CLK _14808_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14739_ hold615/A _14739_/CLK _14739_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08260_ VGND VPWR VGND VPWR _08260_/X _08182_/S _08257_/X _08259_/Y _08280_/B2 sky130_fd_sc_hd__o211a_1
XFILLER_33_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08191_ VGND VPWR VPWR VGND _15519_/D _09792_/A1 _08231_/S hold235/X sky130_fd_sc_hd__mux2_1
X_07211_ VGND VPWR VGND VPWR _08180_/A _07372_/C _07372_/A sky130_fd_sc_hd__xnor2_4
X_07142_ VGND VPWR VGND VPWR _07827_/A _12878_/B _07827_/C _10059_/A _07142_/X sky130_fd_sc_hd__o22a_4
X_07975_ VGND VPWR VGND VPWR _07976_/B _07959_/X _07963_/X _07810_/A _07974_/X sky130_fd_sc_hd__a211o_1
X_09714_ VGND VPWR VPWR VGND _14329_/D fanout24/X _09728_/S hold451/X sky130_fd_sc_hd__mux2_1
XFILLER_27_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09645_ VGND VPWR VPWR VGND _14425_/D hold800/X _09659_/S fanout25/X sky130_fd_sc_hd__mux2_1
XFILLER_43_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09576_ VGND VPWR VPWR VGND _14489_/D hold1001/X _09590_/S fanout24/X sky130_fd_sc_hd__mux2_1
X_08527_ VPWR VGND _15323_/D _08527_/B _11398_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_58_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08458_ VPWR VGND VGND VPWR _08458_/A _08458_/Y _08458_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07409_ VGND VPWR VGND VPWR _07607_/C _07612_/A _07416_/A _07408_/X _10074_/S _07148_/A
+ sky130_fd_sc_hd__a32oi_4
X_13289__406 VPWR VGND VPWR VGND _14564_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_10420_ VGND VPWR VGND VPWR _10420_/X hold773/A _10744_/A2 _10419_/X _10745_/A1 sky130_fd_sc_hd__o211a_1
X_08389_ VGND VPWR VPWR VGND _15388_/D fanout54/X _08405_/S hold610/X sky130_fd_sc_hd__mux2_1
X_10351_ VGND VPWR VPWR VGND _10351_/X hold529/A _10687_/B hold431/A sky130_fd_sc_hd__mux2_1
X_13033__150 VPWR VGND VPWR VGND _14276_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_12917__34 VPWR VGND VPWR VGND _14160_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_14059__1176 VPWR VGND VPWR VGND _15478_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_10282_ VGND VPWR VPWR VGND _10282_/X _10279_/X _10613_/A _10278_/X sky130_fd_sc_hd__mux2_1
X_12021_ VGND VPWR VPWR VGND _12021_/X hold771/A _12190_/S hold227/A sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout560 VPWR VGND _09710_/S _09725_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout593 VPWR VGND _08846_/S _08847_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout582 VPWR VGND _09163_/S _09161_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout571 VPWR VGND _09406_/S _09381_/X VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_8_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_46_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12854_ VGND VPWR VPWR VGND _15578_/D _08132_/Y _12860_/S _09164_/A sky130_fd_sc_hd__mux2_1
X_11805_ VPWR VGND VPWR VGND _11804_/X _12744_/C1 _11803_/X _11805_/Y sky130_fd_sc_hd__a21oi_1
X_15573_ _15573_/Q clkload32/A _15573_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12785_ VPWR VGND VGND VPWR _12789_/A _08080_/Y _10060_/A _12785_/X sky130_fd_sc_hd__o21a_1
X_14524_ hold316/A _14524_/CLK _14524_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11736_ VGND VPWR VPWR VGND _11736_/X _11735_/X _12396_/S _11734_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_41_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11667_ VGND VPWR VGND VPWR _11667_/X _12185_/A1 _11662_/X _11666_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
X_14455_ _14455_/Q _14455_/CLK _14455_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14386_ _14386_/Q clkload9/A _14386_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_10618_ VPWR VGND VGND VPWR _10618_/A _10618_/B _10618_/Y sky130_fd_sc_hd__nor2_1
X_11598_ VGND VPWR VPWR VGND _11598_/X hold956/A _11998_/S hold214/A sky130_fd_sc_hd__mux2_1
X_10549_ VPWR VGND VPWR VGND _10548_/X _10625_/S _10622_/C1 _10549_/X sky130_fd_sc_hd__a21o_1
X_15007_ _15007_/Q _15007_/CLK _15007_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13580__697 VPWR VGND VPWR VGND _14911_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_12219_ VGND VPWR VPWR VGND _12219_/X hold798/A _12219_/S hold722/A sky130_fd_sc_hd__mux2_1
X_07760_ VPWR VGND VGND VPWR _07761_/B _15547_/Q _07760_/B sky130_fd_sc_hd__or2_1
XFILLER_38_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07691_ VGND VPWR VGND VPWR _07691_/X _15129_/Q _15356_/Q _08495_/A2 clone18/X sky130_fd_sc_hd__a22o_4
XFILLER_53_904 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09430_ VGND VPWR VPWR VGND _14622_/D _09443_/S fanout42/X hold1234/X sky130_fd_sc_hd__mux2_4
X_13474__591 VPWR VGND VPWR VGND _14749_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_09361_ VGND VPWR VPWR VGND _14685_/D hold684/X _09376_/S fanout39/X sky130_fd_sc_hd__mux2_1
X_09292_ VGND VPWR VPWR VGND _14749_/D fanout40/X _09304_/S hold508/X sky130_fd_sc_hd__mux2_1
XFILLER_36_1014 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08312_ VGND VPWR VPWR VGND _15507_/D fanout68/X _08318_/S hold1071/X sky130_fd_sc_hd__mux2_1
XANTENNA_23 _14397_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08243_ VPWR VGND VGND VPWR _15448_/Q _07234_/B _08278_/B _08243_/X sky130_fd_sc_hd__o21a_1
XANTENNA_12 _08377_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_45 fanout282/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_1361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_56 _12080_/A2 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_34 _12666_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_13017__134 VPWR VGND VPWR VGND _14260_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_08174_ VPWR VGND VGND VPWR _11284_/B _08174_/Y _08174_/A sky130_fd_sc_hd__nor2_2
XANTENNA_67 _08409_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_89 _14385_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_78 _08366_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07125_ VPWR VGND VPWR VGND _07125_/Y _14834_/Q sky130_fd_sc_hd__inv_2
X_13821__938 VPWR VGND VPWR VGND _15193_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_07958_ VPWR VGND VPWR VGND _07958_/B _07958_/D _07958_/C _07958_/A _07959_/B sky130_fd_sc_hd__or4_1
X_07889_ VPWR VGND VGND VPWR _07993_/A _07889_/B _07890_/D sky130_fd_sc_hd__nor2_1
X_13715__832 VPWR VGND VPWR VGND _15055_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_09628_ _14442_/D fanout91/X fanout87/X _09637_/S _09627_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09559_ _14506_/D fanout94/X fanout90/X _09587_/S _09558_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_15_149 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12570_ VGND VPWR VPWR VGND _12570_/X _14566_/Q _12577_/S _14598_/Q sky130_fd_sc_hd__mux2_1
X_11521_ VGND VPWR VPWR VGND _11521_/X _11520_/X _11537_/S _15471_/Q sky130_fd_sc_hd__mux2_1
X_14240_ _14240_/Q _14240_/CLK _14240_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11452_ VGND VPWR VPWR VGND _11452_/X _11451_/X _11476_/S _15448_/Q sky130_fd_sc_hd__mux2_1
X_10403_ VGND VPWR VGND VPWR _10403_/X _10402_/X _10401_/X _10685_/S _10697_/B1 sky130_fd_sc_hd__a211o_1
X_11383_ VGND VPWR VPWR VGND _11383_/X _14848_/Q _11392_/B _14816_/Q sky130_fd_sc_hd__mux2_1
X_14171_ hold683/A _14171_/CLK _14171_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10334_ VGND VPWR VGND VPWR _10334_/X _10816_/A _10330_/X _10333_/X _11259_/C1 sky130_fd_sc_hd__o211a_1
X_10265_ VPWR VGND _10265_/X _10264_/X _10260_/X _10987_/S _10256_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10196_ VGND VPWR VPWR VGND _10196_/X hold476/A _10567_/S hold484/A sky130_fd_sc_hd__mux2_1
X_12004_ VGND VPWR VGND VPWR _12004_/X _12003_/X _12002_/X _11995_/S _12017_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_78_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout390 VGND VPWR _07872_/Y fanout390/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1023 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_466 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13458__575 VPWR VGND VPWR VGND _14733_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_15625_ _15625_/Q clkload49/A _15625_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12837_ VPWR VGND _12837_/X _15567_/Q _15568_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_12768_ VPWR VGND VGND VPWR _10078_/A _12833_/B _08153_/X _12768_/X sky130_fd_sc_hd__o21a_1
X_15556_ _15556_/Q clkload44/A _15556_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15487_ hold782/A _15487_/CLK _15487_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12699_ VPWR VGND VGND VPWR _12699_/X hold329/A _12708_/S sky130_fd_sc_hd__or2_1
X_11719_ VGND VPWR VPWR VGND _11719_/X hold804/A _11748_/S hold461/A sky130_fd_sc_hd__mux2_1
X_14507_ hold214/A _14507_/CLK _14507_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14438_ _14438_/Q _14438_/CLK _14438_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold805 hold805/X hold805/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 hold827/X hold827/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 hold816/X hold816/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ hold843/A _14369_/CLK _14369_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold838 hold838/X hold838/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 hold849/X hold849/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08930_ VPWR VGND VPWR VGND _09885_/C hold212/A _09970_/B _14148_/Q _14147_/Q sky130_fd_sc_hd__or4b_2
XFILLER_48_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08861_ VPWR VGND VPWR VGND hold819/A _09900_/A _14142_/Q _08862_/C sky130_fd_sc_hd__or3_1
X_07812_ VPWR VGND _07813_/B _07897_/A _07812_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_57_539 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08792_ VGND VPWR VPWR VGND _15217_/D _08811_/S clone46/A hold1150/X sky130_fd_sc_hd__mux2_4
X_07743_ _08076_/A _07741_/X _07743_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_65_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07674_ VGND VPWR VPWR VGND _15539_/D fanout68/X _08231_/S hold306/X sky130_fd_sc_hd__mux2_1
X_14058__1175 VPWR VGND VPWR VGND _15477_/CLK clkload29/A sky130_fd_sc_hd__inv_2
XFILLER_77_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09413_ VGND VPWR VPWR VGND _14636_/D hold460/X _09414_/S fanout98/X sky130_fd_sc_hd__mux2_1
XFILLER_80_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_55_1445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_1418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09344_ VGND VPWR VPWR VGND _14700_/D hold648/X _09345_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
X_09275_ VGND VPWR VPWR VGND _14768_/D fanout97/X _09275_/S hold611/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13251__368 VPWR VGND VPWR VGND _14526_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_08226_ VPWR VGND VGND VPWR _15449_/Q _12845_/A _08278_/B _08226_/X sky130_fd_sc_hd__o21a_1
X_08157_ VPWR VGND VGND VPWR _08240_/A _08157_/Y _08157_/B sky130_fd_sc_hd__nand2_1
X_07108_ VPWR VGND VPWR VGND _07108_/Y _14828_/Q sky130_fd_sc_hd__inv_2
X_08088_ VGND VPWR VGND VPWR _08088_/X _08083_/A _08066_/B _08085_/X _08087_/Y sky130_fd_sc_hd__o211a_1
X_10050_ VPWR VGND _15636_/D _10050_/B _10051_/B VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_75_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_57_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13145__262 VPWR VGND VPWR VGND _14420_/CLK clkload17/A sky130_fd_sc_hd__inv_2
XFILLER_44_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10952_ VGND VPWR VPWR VGND _10952_/X hold774/A _11179_/S hold991/A sky130_fd_sc_hd__mux2_1
X_10883_ VPWR VGND VPWR VGND _10880_/X _10890_/A _10882_/X _10883_/X sky130_fd_sc_hd__a21o_1
X_15410_ hold361/A _15410_/CLK _15410_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12622_ VGND VPWR VPWR VGND _12622_/X hold941/A _12635_/B hold487/A sky130_fd_sc_hd__mux2_1
X_15341_ _15341_/Q _15341_/CLK _15341_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12553_ VGND VPWR VPWR VGND _12553_/X hold783/A _12664_/S hold708/A sky130_fd_sc_hd__mux2_1
X_11504_ VGND VPWR VPWR VGND _15085_/D _11503_/X _11538_/S hold1332/X sky130_fd_sc_hd__mux2_1
X_15272_ _15272_/Q _15272_/CLK _15272_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13843__960 VPWR VGND VPWR VGND _15215_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_14223_ hold347/A _14223_/CLK _14223_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12484_ VGND VPWR VGND VPWR _12484_/X _15505_/Q _12488_/A2 _12470_/S _12483_/X sky130_fd_sc_hd__o211a_1
X_11435_ VGND VPWR VGND VPWR _14932_/D hold1434/X _11439_/A2 _11434_/X _09977_/A sky130_fd_sc_hd__o211a_1
XFILLER_32_1286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14154_ _14154_/Q _14154_/CLK input1/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11366_ VPWR VGND VGND VPWR _11368_/A _11368_/B _11418_/S sky130_fd_sc_hd__nor2_1
X_10317_ VPWR VGND VGND VPWR _10317_/X hold152/A _11098_/S sky130_fd_sc_hd__or2_1
X_11297_ VGND VPWR VPWR VGND _11298_/B _14817_/Q _11299_/S _14385_/Q sky130_fd_sc_hd__mux2_1
X_10248_ VPWR VGND VGND VPWR _11210_/A _10248_/B _10248_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_78_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10179_ VPWR VGND VPWR VGND _10178_/X _10677_/S _10697_/B1 _10179_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_1079 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14987_ hold757/A _14987_/CLK _14987_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_745 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15608_ _15608_/Q clkload27/A _15608_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07390_ VPWR VGND VPWR VGND _08007_/A _07982_/B _07389_/Y _07397_/B sky130_fd_sc_hd__a21oi_1
X_15539_ hold306/A _15539_/CLK _15539_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09060_ VPWR VGND VGND VPWR _09764_/A _15639_/Q _09557_/A sky130_fd_sc_hd__nand2_2
X_08011_ VPWR VGND VPWR VGND _10074_/A0 _07264_/B _10074_/A1 _08011_/X _07262_/X sky130_fd_sc_hd__a22o_1
X_13088__205 VPWR VGND VPWR VGND _14331_/CLK clkload21/A sky130_fd_sc_hd__inv_2
Xhold602 hold602/X hold602/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 hold613/X hold613/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 hold635/X hold635/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 hold624/X hold624/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 hold679/X hold679/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ VPWR VGND VPWR VGND _15568_/Q _15567_/Q _15569_/Q _12842_/B sky130_fd_sc_hd__or3_1
Xhold668 hold668/X hold668/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 hold646/X hold646/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 hold657/X hold657/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ VGND VPWR VGND VPWR _15136_/D hold1277/X _08919_/A2 _08912_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
X_13129__246 VPWR VGND VPWR VGND _14372_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_09893_ VPWR VGND VGND VPWR _09893_/A _09907_/S _09893_/Y sky130_fd_sc_hd__nor2_1
Xhold1313 hold1313/X _15140_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1302 hold1302/X _15345_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08844_ VGND VPWR VPWR VGND _15169_/D _09792_/A1 _08844_/S hold797/X sky130_fd_sc_hd__mux2_1
Xhold1324 _10021_/A _15624_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 hold1335/X _14850_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 _10037_/A _15631_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1357 hold1357/X _14730_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 _09278_/A _14762_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08775_ VGND VPWR VPWR VGND _15231_/D _09863_/A0 _08776_/S hold267/X sky130_fd_sc_hd__mux2_1
Xhold1379 hold1379/X _14136_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07726_ VPWR VGND VPWR VGND _07827_/D _15586_/Q _07714_/X _07728_/B sky130_fd_sc_hd__a21o_1
X_13786__903 VPWR VGND VPWR VGND _15158_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_07657_ VGND VPWR VGND VPWR _10074_/A1 _07653_/A _07859_/B _07657_/X _07167_/Y sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07588_ VPWR VGND VPWR VGND _07588_/X _07125_/Y _09007_/B _07586_/C _07126_/Y _11284_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_25_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09327_ VGND VPWR VPWR VGND _14717_/D hold742/X _09327_/S fanout39/X sky130_fd_sc_hd__mux2_1
Xclone13 VGND VPWR clone13/X clone13/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_13827__944 VPWR VGND VPWR VGND _15199_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_09258_ VGND VPWR VPWR VGND _14785_/D fanout35/X _09268_/S hold749/X sky130_fd_sc_hd__mux2_1
Xclone46 VPWR VGND clone46/X clone46/A VPWR VGND sky130_fd_sc_hd__buf_6
X_09189_ VGND VPWR VPWR VGND _14902_/D hold344/X _09197_/S _09825_/A1 sky130_fd_sc_hd__mux2_1
X_08209_ VGND VPWR VGND VPWR _15611_/Q _08220_/A _08208_/X _08209_/X _08299_/A2 sky130_fd_sc_hd__a2bb2o_1
X_11220_ VPWR VGND VGND VPWR _11220_/X hold210/A _11223_/S sky130_fd_sc_hd__or2_1
XFILLER_68_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11151_ VGND VPWR VGND VPWR _11151_/X _15027_/Q _11252_/A2 _11150_/X _11143_/S sky130_fd_sc_hd__o211a_1
X_10102_ VGND VPWR VPWR VGND _10102_/X hold851/A _10609_/S hold531/A sky130_fd_sc_hd__mux2_1
X_11082_ VGND VPWR VPWR VGND _11082_/X _14630_/Q _11091_/S _14662_/Q sky130_fd_sc_hd__mux2_1
X_10033_ VPWR VGND VGND VPWR _10035_/B _10033_/B _15629_/D sky130_fd_sc_hd__nor2_1
X_14910_ hold337/A _14910_/CLK _14910_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_7_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14841_ _14841_/Q clkload28/A _14841_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_1173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_542 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11984_ VGND VPWR VPWR VGND _11984_/X hold459/A _11998_/S hold410/A sky130_fd_sc_hd__mux2_1
X_14772_ hold753/A _14772_/CLK _14772_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10935_ VGND VPWR VPWR VGND _10935_/X hold787/A _11179_/S hold825/A sky130_fd_sc_hd__mux2_1
X_10866_ VGND VPWR VGND VPWR _10866_/X _10865_/X _10864_/X _11110_/A _12868_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_32_726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12605_ VGND VPWR VPWR VGND _12605_/X hold751/A _12623_/S hold643/A sky130_fd_sc_hd__mux2_1
X_15324_ _15324_/Q _15324_/CLK _15324_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10797_ VGND VPWR VPWR VGND _10797_/X hold438/A _11204_/S hold268/A sky130_fd_sc_hd__mux2_1
X_13273__390 VPWR VGND VPWR VGND _14548_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_12536_ VGND VPWR VPWR VGND _12536_/X _12533_/X _12536_/S _12532_/X sky130_fd_sc_hd__mux2_1
X_12467_ VGND VPWR VPWR VGND _12467_/X hold597/A _12479_/S hold413/A sky130_fd_sc_hd__mux2_1
X_15255_ hold348/A _15255_/CLK _15255_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11418_ VGND VPWR VPWR VGND _11418_/X _11356_/X _11418_/S _15702_/A sky130_fd_sc_hd__mux2_1
X_14206_ _14206_/Q _14206_/CLK _14206_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15186_ hold772/A _15186_/CLK _15186_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14137_ _14137_/Q _14137_/CLK _14137_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12398_ VGND VPWR VPWR VGND _12399_/B _12397_/Y _12472_/S _12389_/Y sky130_fd_sc_hd__mux2_1
X_11349_ VGND VPWR VPWR VGND _11349_/X _14927_/Q _11355_/S hold1224/X sky130_fd_sc_hd__mux2_1
X_14057__1174 VPWR VGND VPWR VGND _15429_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_80_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13620__737 VPWR VGND VPWR VGND _14960_/CLK clkload38/A sky130_fd_sc_hd__inv_2
XFILLER_80_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1308 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_78_1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08560_ VPWR VGND VGND VPWR _08559_/A _08559_/B _07534_/B _08560_/X sky130_fd_sc_hd__o21a_1
X_08491_ VPWR VGND _08491_/X _11302_/B _08491_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07511_ VPWR VGND VGND VPWR _07512_/B _15465_/Q _07511_/B sky130_fd_sc_hd__or2_1
XFILLER_78_1297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07442_ VPWR VGND VGND VPWR _08545_/A _15458_/Q _07714_/A sky130_fd_sc_hd__or2_1
X_13514__631 VPWR VGND VPWR VGND _14789_/CLK clkload46/A sky130_fd_sc_hd__inv_2
Xfanout29 VGND VPWR _08014_/X fanout29/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07373_ _08137_/C _08162_/A _08180_/A _08180_/B _07371_/X _07372_/X VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__o311a_1
X_09112_ VGND VPWR VPWR VGND _14983_/D hold419/X _09128_/S fanout34/X sky130_fd_sc_hd__mux2_1
X_09043_ VGND VPWR VPWR VGND _15047_/D hold420/X _09051_/S fanout33/X sky130_fd_sc_hd__mux2_1
Xhold410 hold410/X hold410/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 hold432/X hold432/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 hold443/X hold443/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold421 hold421/X hold421/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 hold454/X hold454/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 hold476/X hold476/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 hold487/X hold487/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 hold465/X hold465/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ VGND VPWR _09947_/C _09945_/Y _14129_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold498 hold498/X hold498/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09876_ VPWR VGND VPWR VGND _09875_/Y _09878_/B _09882_/A _14151_/D sky130_fd_sc_hd__a21oi_1
Xhold1132 hold1132/X _14726_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 hold1121/X _15058_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_645 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1110 hold1110/X _15024_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Left_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08827_ VGND VPWR VPWR VGND _15186_/D fanout56/X _08846_/S hold772/X sky130_fd_sc_hd__mux2_1
Xhold1143 hold1143/X _14142_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 hold1154/X _14246_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 hold1176/X _15344_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_678 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1165 hold1165/X _14504_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 hold1187/X _14840_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1198 hold1198/X _15335_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ VGND VPWR VPWR VGND _15248_/D clone100/X _08776_/S hold630/X sky130_fd_sc_hd__mux2_1
X_07709_ VPWR VGND VGND VPWR _07710_/B _15564_/Q _07709_/B sky130_fd_sc_hd__or2_1
X_08689_ VGND VPWR VGND VPWR _15285_/D hold1295/X _08701_/A2 _08688_/X _12085_/C1
+ sky130_fd_sc_hd__o211a_1
X_10720_ VGND VPWR VPWR VGND _10724_/B hold749/A _10720_/S hold334/A sky130_fd_sc_hd__mux2_1
XFILLER_13_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13257__374 VPWR VGND VPWR VGND _14532_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_10651_ VGND VPWR VGND VPWR _10651_/X _10557_/A _10647_/X _10650_/X _10717_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_10_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10582_ VPWR VGND VGND VPWR _10582_/X hold437/A _10730_/S sky130_fd_sc_hd__or2_1
X_12321_ VGND VPWR VGND VPWR _12321_/X _12580_/A1 _12317_/X _12320_/X _12572_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_16_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12252_ VGND VPWR VPWR VGND _12252_/X hold947/A _12578_/S hold684/A sky130_fd_sc_hd__mux2_1
X_15040_ hold696/A _15040_/CLK _15040_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11203_ VGND VPWR VPWR VGND _11203_/X _14217_/Q _11204_/S hold222/A sky130_fd_sc_hd__mux2_1
X_12962__79 VPWR VGND VPWR VGND _14205_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_12183_ VGND VPWR VPWR VGND _12183_/X _14878_/Q _12183_/S hold380/A sky130_fd_sc_hd__mux2_1
X_11134_ VPWR VGND VPWR VGND _11133_/X _11245_/A1 _11132_/X _11134_/Y sky130_fd_sc_hd__a21oi_1
X_11065_ VGND VPWR VPWR VGND _11065_/X _11064_/X _11176_/S _11063_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10016_ VGND VPWR VPWR VGND _10016_/A _15622_/D _10017_/C sky130_fd_sc_hd__xor2_1
XFILLER_7_1257 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_48_177 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_37_829 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_818 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14824_ _14824_/Q clkload28/A _14824_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11967_ VPWR VGND VGND VPWR _11968_/S _11963_/X _12184_/C1 _11967_/X sky130_fd_sc_hd__o21a_1
X_14755_ hold413/A _14755_/CLK _14755_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10918_ VGND VPWR VGND VPWR _10918_/X _10917_/X _10916_/X _11235_/A1 _10918_/C1 sky130_fd_sc_hd__a211o_1
X_11898_ VPWR VGND VGND VPWR _11879_/X _11896_/X _07913_/Y _11897_/X _11898_/X sky130_fd_sc_hd__o22a_1
X_14686_ _14686_/Q _14686_/CLK _14686_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10849_ VGND VPWR VPWR VGND _10853_/B hold963/A _10850_/S hold228/A sky130_fd_sc_hd__mux2_1
X_15307_ _15307_/Q _15307_/CLK _15307_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12519_ VGND VPWR VPWR VGND _12519_/X hold627/A _12671_/S hold272/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15238_ hold232/A _15238_/CLK _15238_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13050__167 VPWR VGND VPWR VGND _14293_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_15169_ hold797/A _15169_/CLK _15169_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout208 VPWR VGND _12375_/S _07978_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_07991_ VGND VPWR VPWR VGND _07991_/X _07974_/B1 _07987_/X _07886_/A _07990_/X sky130_fd_sc_hd__o2bb2a_1
Xfanout219 VPWR VGND _12017_/C1 _12115_/C1 VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_80_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09730_ VPWR VGND VPWR VGND _09730_/Y _09757_/S sky130_fd_sc_hd__inv_2
XFILLER_67_420 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xtt_um_femto_902 uio_out[5] tt_um_femto_902/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09661_ VPWR VGND VGND VPWR hold1378/X _09687_/S _09661_/Y sky130_fd_sc_hd__nand2b_1
X_08612_ VGND VPWR VGND VPWR _08612_/X _08582_/A _08615_/B1 hold1054/X _08611_/Y sky130_fd_sc_hd__a211o_1
XFILLER_55_648 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_136 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09592_ VPWR VGND VPWR VGND _09592_/Y _09622_/S sky130_fd_sc_hd__inv_2
X_08543_ VPWR VGND VGND VPWR _08566_/A _08566_/B _08544_/B sky130_fd_sc_hd__nor2_1
X_08474_ VPWR VGND VGND VPWR _08474_/X _15339_/Q _08482_/B sky130_fd_sc_hd__or2_1
XFILLER_56_1392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07425_ _07425_/X _12878_/A _07703_/A _07827_/B _07807_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_51_887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07356_ VPWR VGND VPWR VGND _07355_/Y _08083_/A _07354_/X _07356_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_1207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07287_ VPWR VGND VGND VPWR _07288_/A _07946_/A _07287_/Y sky130_fd_sc_hd__nor2_1
X_09026_ VPWR VGND VPWR VGND _09026_/X _09799_/A _09095_/B sky130_fd_sc_hd__or2_2
XFILLER_3_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold251 hold251/X hold251/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/X hold240/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/X hold262/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/X hold295/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/X hold273/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/X hold284/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ VGND VPWR _09931_/C _09928_/Y _14134_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
Xfanout742 VPWR VGND _08220_/A _07828_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout731 VGND VPWR _12751_/A2 _12677_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout720 VGND VPWR _12195_/B1 _12047_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout753 VPWR VGND _12817_/A _12790_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout764 VGND VPWR _08002_/A2 _07929_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout775 VGND VPWR _07414_/Y _08280_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout797 VPWR VGND _08626_/A fanout802/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout786 VPWR VGND _11340_/A _09938_/A VPWR VGND sky130_fd_sc_hd__buf_4
X_09859_ VGND VPWR VPWR VGND _14163_/D hold506/X _09867_/S _09859_/A0 sky130_fd_sc_hd__mux2_1
X_12870_ VGND VPWR VPWR VGND _15594_/D _11210_/A _12870_/S _15594_/Q sky130_fd_sc_hd__mux2_1
X_11821_ VPWR VGND VGND VPWR _11821_/X hold759/A _12372_/S sky130_fd_sc_hd__or2_1
XANTENNA_113 _09825_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_102 _10705_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_14540_ hold647/A _14540_/CLK _14540_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14056__1173 VPWR VGND VPWR VGND _15428_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_11752_ VPWR VGND VGND VPWR _11733_/Y _11751_/X _12380_/B _15449_/Q _15449_/D _12492_/C1
+ sky130_fd_sc_hd__o221a_1
X_10703_ VPWR VGND VGND VPWR _10703_/X _10703_/A _10703_/B sky130_fd_sc_hd__or2_1
X_14471_ hold582/A _14471_/CLK _14471_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11683_ VPWR VGND VGND VPWR _11683_/X _12476_/S _11683_/B sky130_fd_sc_hd__or2_1
X_10634_ VGND VPWR VGND VPWR _10634_/X _10631_/X _10633_/X _10634_/A1 _10634_/C1 sky130_fd_sc_hd__a211o_1
X_12304_ VGND VPWR VGND VPWR _12304_/X _12303_/X _12302_/X _12748_/A1 _12748_/C1 sky130_fd_sc_hd__a211o_1
X_10565_ VGND VPWR VPWR VGND _10565_/X hold906/A _10735_/S hold820/A sky130_fd_sc_hd__mux2_1
X_10496_ VGND VPWR VPWR VGND _10496_/X _10493_/X _10510_/S _10492_/X sky130_fd_sc_hd__mux2_1
X_12235_ VPWR VGND VGND VPWR _12235_/X hold855/A _12578_/S sky130_fd_sc_hd__or2_1
X_15023_ _15023_/Q _15023_/CLK _15023_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12166_ VGND VPWR VPWR VGND _12166_/X _12163_/X _12174_/S _12162_/X sky130_fd_sc_hd__mux2_1
X_11117_ VPWR VGND VGND VPWR _11117_/X _14406_/Q _11117_/B sky130_fd_sc_hd__or2_1
XFILLER_42_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13691__808 VPWR VGND VPWR VGND _15031_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_12097_ VGND VPWR VPWR VGND _12097_/X _14457_/Q _12097_/S _14745_/Q sky130_fd_sc_hd__mux2_1
XFILLER_77_762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11048_ VGND VPWR VPWR VGND _11048_/X hold695/A _11054_/S hold389/A sky130_fd_sc_hd__mux2_1
X_14807_ _14807_/Q _14807_/CLK _14807_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13732__849 VPWR VGND VPWR VGND _15104_/CLK clkload30/A sky130_fd_sc_hd__inv_2
XFILLER_64_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_45_681 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_75_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14738_ hold282/A _14738_/CLK _14738_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14669_ hold477/A _14669_/CLK _14669_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08190_ VGND VPWR VGND VPWR _08249_/A2 _15612_/Q _08189_/Y _08190_/X _08178_/X sky130_fd_sc_hd__a211o_4
X_07210_ VPWR VGND VGND VPWR _07210_/X _15451_/Q _07372_/C sky130_fd_sc_hd__or2_1
X_13585__702 VPWR VGND VPWR VGND _14916_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_07141_ VGND VPWR VGND VPWR _12878_/B _07703_/A _15574_/Q _15572_/Q _07141_/A sky130_fd_sc_hd__or4b_4
XFILLER_12_1240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13626__743 VPWR VGND VPWR VGND _14966_/CLK clkload33/A sky130_fd_sc_hd__inv_2
XFILLER_10_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07974_ _07974_/X _07970_/X _07971_/Y _07973_/X _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09713_ VGND VPWR VPWR VGND _14330_/D fanout29/X _09721_/S hold700/X sky130_fd_sc_hd__mux2_1
XFILLER_55_423 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09644_ VGND VPWR VPWR VGND _14426_/D hold874/X _09657_/S fanout29/X sky130_fd_sc_hd__mux2_1
XFILLER_35_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09575_ VGND VPWR VPWR VGND _14490_/D hold996/X _09588_/S fanout29/X sky130_fd_sc_hd__mux2_1
X_08526_ VPWR VGND VPWR VGND _08534_/B1 _15322_/Q _08503_/A _08527_/B hold1392/X sky130_fd_sc_hd__a22o_1
XFILLER_58_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08457_ VGND VPWR VGND VPWR _15348_/D hold1344/X _08458_/B _08456_/X _11308_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_19_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_695 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07408_ VGND VPWR VGND VPWR _07408_/X _07607_/B _07410_/B _07612_/A _07411_/A sky130_fd_sc_hd__a211o_1
X_08388_ VGND VPWR VPWR VGND _15389_/D clone55/A _08405_/S hold687/X sky130_fd_sc_hd__mux2_1
X_07339_ VPWR VGND VPWR VGND _07665_/A _07668_/A _07339_/B sky130_fd_sc_hd__or2_2
X_10350_ VGND VPWR VPWR VGND _10354_/B hold485/A _10687_/B hold213/A sky130_fd_sc_hd__mux2_1
X_13369__486 VPWR VGND VPWR VGND _14644_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_09009_ VGND VPWR VGND VPWR hold972/A hold971/X _09015_/A2 _09008_/X _11327_/A sky130_fd_sc_hd__o211a_1
X_10281_ VGND VPWR VGND VPWR _10281_/X _10614_/A1 _10277_/X _10280_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
X_12020_ VGND VPWR VPWR VGND _12024_/B hold854/A _12190_/S hold175/A sky130_fd_sc_hd__mux2_1
X_12932__49 VPWR VGND VPWR VGND _14175_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
Xfanout550 VPWR VGND _07567_/B clone13/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout572 VPWR VGND _09408_/S _09411_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout561 _09725_/S _09694_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout583 VPWR VGND _09161_/S _09129_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout594 VPWR VGND _08844_/S _08847_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_12853_ VGND VPWR VPWR VGND _15577_/D _07591_/Y _12860_/S _15577_/Q sky130_fd_sc_hd__mux2_1
X_11804_ VGND VPWR VPWR VGND _11804_/X _11801_/X _12591_/S _11800_/X sky130_fd_sc_hd__mux2_1
X_12784_ VGND VPWR VPWR VGND _15553_/D _12783_/Y _12782_/X _12807_/A1 _12807_/B1 _15553_/Q
+ sky130_fd_sc_hd__a32o_1
X_15572_ _15572_/Q clkload27/A _15572_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_38_Left_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_72_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14523_ hold291/A _14523_/CLK _14523_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_342 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11735_ VGND VPWR VPWR VGND _11735_/X _14351_/Q _12409_/B hold675/A sky130_fd_sc_hd__mux2_1
XFILLER_15_887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_30_846 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14454_ hold631/A _14454_/CLK _14454_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11666_ VGND VPWR VGND VPWR _11666_/X _11665_/X _11664_/X _11948_/S _12184_/C1 sky130_fd_sc_hd__a211o_1
X_13313__430 VPWR VGND VPWR VGND _14588_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_14385_ VGND VPWR VGND VPWR _14385_/Q _14385_/D clkload55/A sky130_fd_sc_hd__dfxtp_4
X_11597_ VGND VPWR VGND VPWR _11597_/X _11594_/X _11596_/X _12099_/A1 _12101_/A1 sky130_fd_sc_hd__a211o_1
X_10617_ VGND VPWR VPWR VGND _10618_/B _10616_/Y _10617_/S _10608_/Y sky130_fd_sc_hd__mux2_1
X_10548_ VGND VPWR VPWR VGND _10548_/X _14874_/Q _10627_/S hold361/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_47_Left_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10479_ VGND VPWR VPWR VGND _10479_/X hold718/A _10479_/S hold248/A sky130_fd_sc_hd__mux2_1
X_15006_ _15006_/Q _15006_/CLK _15006_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12218_ VGND VPWR VGND VPWR _12218_/X _12217_/X _12216_/X _12230_/A1 _12226_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_9_1116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12149_ VGND VPWR VPWR VGND _12149_/X hold393/A _12149_/S hold660/A sky130_fd_sc_hd__mux2_1
X_13162__279 VPWR VGND VPWR VGND _14437_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_07690_ VGND VPWR VGND VPWR _15356_/Q _08495_/A2 _15129_/Q _07690_/Y _07873_/B1 sky130_fd_sc_hd__a22oi_4
XFILLER_25_607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_80_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09360_ VGND VPWR VPWR VGND _14686_/D _09376_/S hold1185/X clone44/X sky130_fd_sc_hd__mux2_4
X_08311_ VGND VPWR VPWR VGND _15508_/D _08332_/S clone111/X hold1267/X sky130_fd_sc_hd__mux2_4
X_09291_ VGND VPWR VPWR VGND _14750_/D clone6/X _09307_/S hold620/X sky130_fd_sc_hd__mux2_1
XFILLER_75_1097 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08242_ VGND VPWR VGND VPWR _08242_/X _08277_/S _08241_/X _08240_/Y _08280_/B2 sky130_fd_sc_hd__o211a_1
XANTENNA_13 _08745_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_46 fanout382/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_57 _12080_/A2 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_13056__173 VPWR VGND VPWR VGND _14299_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XANTENNA_24 _14397_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_35 _12666_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_79 _08372_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08173_ VGND VPWR VPWR VGND _08214_/A _08173_/Y _07331_/A _08195_/A sky130_fd_sc_hd__o21ai_4
XANTENNA_68 _08409_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07124_ VPWR VGND VPWR VGND _11367_/D _14853_/Q sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_65_Left_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13860__977 VPWR VGND VPWR VGND _15232_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
XFILLER_47_1133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_47_1177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14055__1172 VPWR VGND VPWR VGND _15427_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XFILLER_60_1333 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07957_ VPWR VGND VPWR VGND _08270_/A1 _07331_/A _07598_/Y _07976_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13754__871 VPWR VGND VPWR VGND _15126_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_07888_ VGND VPWR _07888_/B _07889_/B _07888_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_56_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09627_ VPWR VGND VGND VPWR hold1385/X _09637_/S _09627_/Y sky130_fd_sc_hd__nand2b_1
X_09558_ VPWR VGND _09558_/X _09834_/B _09486_/B _09164_/A _14506_/Q VGND VPWR sky130_fd_sc_hd__a31o_1
X_08509_ VPWR VGND VPWR VGND _08534_/B1 _15330_/Q _08503_/A _08510_/B hold1437/X sky130_fd_sc_hd__a22o_1
XFILLER_62_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11520_ VGND VPWR VPWR VGND _11520_/X _15092_/Q _11529_/S _15090_/Q sky130_fd_sc_hd__mux2_1
X_09489_ _14570_/D fanout94/X fanout90/X _09487_/Y _09488_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_24_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_23_194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11451_ VGND VPWR VPWR VGND _11451_/X _15069_/Q _11475_/S _15067_/Q sky130_fd_sc_hd__mux2_1
X_10402_ VGND VPWR VPWR VGND _10402_/X hold910/A _10696_/S hold725/A sky130_fd_sc_hd__mux2_1
X_11382_ VGND VPWR VPWR VGND _14847_/D _11381_/X _11382_/S hold1306/X sky130_fd_sc_hd__mux2_1
X_14170_ hold533/A _14170_/CLK _14170_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10333_ VPWR VGND VGND VPWR _10333_/X _10333_/A _10333_/B sky130_fd_sc_hd__or2_1
X_10264_ VGND VPWR VGND VPWR _10264_/X _10261_/X _10263_/X _11235_/A1 _10930_/C1 sky130_fd_sc_hd__a211o_1
X_10195_ VGND VPWR VPWR VGND _10195_/X hold863/A _10972_/S hold439/A sky130_fd_sc_hd__mux2_1
X_12003_ VGND VPWR VPWR VGND _12003_/X hold669/A _12005_/S hold236/A sky130_fd_sc_hd__mux2_1
Xfanout380 VGND VPWR fanout381/X _11205_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout391 VGND VPWR _10593_/A1 _10557_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_15624_ _15624_/Q clkload49/A _15624_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12836_ VGND VPWR VGND VPWR _15567_/D _08290_/B _11476_/S _11477_/S _07082_/Y sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_1_Left_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15555_ _15555_/Q clkload27/A _15555_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14506_ _14506_/Q _14506_/CLK _14506_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12767_ VGND VPWR VPWR VGND _15549_/D _12766_/X _12765_/Y _12834_/C1 _12807_/B1 _15549_/Q
+ sky130_fd_sc_hd__a32o_1
X_12698_ VGND VPWR VPWR VGND _12698_/X _12697_/X _12698_/S _12696_/X sky130_fd_sc_hd__mux2_1
X_11718_ VGND VPWR VPWR VGND _11718_/X hold664/A _11748_/S hold267/A sky130_fd_sc_hd__mux2_1
X_15486_ hold958/A _15486_/CLK _15486_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11649_ VPWR VGND VPWR VGND _11648_/X _12185_/A1 _11647_/X _11649_/Y sky130_fd_sc_hd__a21oi_1
X_14437_ _14437_/Q _14437_/CLK _14437_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14368_ _14368_/Q _14368_/CLK _14368_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold817 hold817/X hold817/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold806 hold806/X hold806/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 hold828/X hold828/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14299_ hold196/A _14299_/CLK _14299_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold839 hold839/X hold839/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13697__814 VPWR VGND VPWR VGND _15037_/CLK clkload49/A sky130_fd_sc_hd__inv_2
XFILLER_48_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08860_ VPWR VGND VGND VPWR _14142_/Q _09900_/A _08860_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07811_ VPWR VGND VPWR VGND _07811_/B _07899_/A _07811_/A _07897_/A sky130_fd_sc_hd__or3_1
X_13738__855 VPWR VGND VPWR VGND _15110_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_08791_ VGND VPWR VPWR VGND _15218_/D fanout58/X _08808_/S hold174/X sky130_fd_sc_hd__mux2_1
X_07742_ VPWR VGND VGND VPWR _07743_/B _15554_/Q _07742_/B sky130_fd_sc_hd__or2_1
X_07673_ VPWR VGND VGND VPWR _07673_/X _07673_/A _07673_/B sky130_fd_sc_hd__or2_1
X_09412_ VGND VPWR VPWR VGND _14637_/D hold333/X _09414_/S _09865_/A0 sky130_fd_sc_hd__mux2_1
X_09343_ VGND VPWR VPWR VGND _14701_/D hold401/X _09345_/S _09691_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_61_790 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_55_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09274_ VGND VPWR VPWR VGND _14769_/D fanout98/X _09275_/S hold427/X sky130_fd_sc_hd__mux2_1
X_08225_ VGND VPWR VGND VPWR _08225_/X _08182_/S _08222_/X _08224_/X _08225_/C1 sky130_fd_sc_hd__o211a_1
X_08156_ VGND VPWR _08156_/B _08157_/B _08162_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07107_ VPWR VGND VPWR VGND _07107_/Y _14832_/Q sky130_fd_sc_hd__inv_2
X_13892__1009 VPWR VGND VPWR VGND _15264_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
XFILLER_49_1228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08087_ VPWR VGND VPWR VGND _11440_/B _15076_/Q _08086_/X _08087_/Y sky130_fd_sc_hd__a21oi_1
X_12902__19 VPWR VGND VPWR VGND _14144_/CLK clkload29/A sky130_fd_sc_hd__inv_2
XFILLER_57_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08989_ VPWR VGND VGND VPWR _09873_/A _08989_/B _08989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13490__607 VPWR VGND VPWR VGND _14765_/CLK clkload26/A sky130_fd_sc_hd__inv_2
XFILLER_44_713 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10951_ VPWR VGND VGND VPWR _11173_/A _10951_/B _10951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10882_ VPWR VGND VPWR VGND _10881_/X _11110_/A _12868_/A1 _10882_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12621_ VPWR VGND VGND VPWR _12658_/A _12621_/B _12621_/Y sky130_fd_sc_hd__nor2_1
X_13531__648 VPWR VGND VPWR VGND _14862_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_15340_ _15340_/Q _15340_/CLK _15340_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12552_ VGND VPWR VPWR VGND _12552_/X _14437_/Q _12664_/S hold436/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11503_ VGND VPWR VPWR VGND _11503_/X _11502_/X _11537_/S _15465_/Q sky130_fd_sc_hd__mux2_1
X_15271_ hold976/A _15271_/CLK _15271_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12483_ VPWR VGND VGND VPWR _12483_/X hold179/A _12716_/S sky130_fd_sc_hd__or2_1
X_11434_ VGND VPWR VGND VPWR _11434_/X _14932_/Q _07109_/Y _11439_/A2 sky130_fd_sc_hd__a21bo_1
X_14222_ hold253/A _14222_/CLK _14222_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13384__501 VPWR VGND VPWR VGND _14659_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_11365_ VGND VPWR _11367_/D _14851_/Q _11368_/B _14852_/Q _14854_/Q VPWR VGND sky130_fd_sc_hd__and4b_1
X_14153_ _14153_/Q clkload43/A _14153_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10316_ VGND VPWR VPWR VGND _10316_/X hold605/A _11098_/S hold308/A sky130_fd_sc_hd__mux2_1
X_11296_ VPWR VGND _14816_/D _11296_/B _11296_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_4_864 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10247_ VGND VPWR VPWR VGND _10248_/B _10246_/Y _10987_/S _10238_/Y sky130_fd_sc_hd__mux2_1
X_13425__542 VPWR VGND VPWR VGND _14700_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_10178_ VGND VPWR VPWR VGND _10178_/X hold927/A _10484_/B hold445/A sky130_fd_sc_hd__mux2_1
X_14986_ hold891/A _14986_/CLK _14986_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_724 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_510 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12819_ VPWR VGND VGND VPWR _12818_/X _12834_/C1 _07527_/X _12817_/Y _15562_/D sky130_fd_sc_hd__o22a_1
XFILLER_50_738 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15607_ _15607_/Q clkload27/A _15607_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_481 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15538_ hold272/A _15538_/CLK _15538_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14054__1171 VPWR VGND VPWR VGND _15426_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_15469_ _15469_/Q clkload36/A _15469_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08010_ VPWR VGND VGND VPWR _08010_/X _08010_/A _08066_/B sky130_fd_sc_hd__or2_1
X_12968__85 VPWR VGND VPWR VGND _14211_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
Xhold603 hold603/X hold603/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 hold636/X hold636/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 hold625/X hold625/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 hold614/X hold614/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 hold658/X hold658/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ VPWR VGND VGND VPWR _15568_/Q _15567_/Q _09961_/Y sky130_fd_sc_hd__nor2_1
Xhold647 hold647/X hold647/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 hold669/X hold669/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ VPWR VGND VGND VPWR _08912_/X _15136_/Q _08926_/B sky130_fd_sc_hd__or2_1
X_13168__285 VPWR VGND VPWR VGND _14443_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_09892_ VPWR VGND VPWR VGND _15477_/D _09892_/C _09892_/A _09907_/S sky130_fd_sc_hd__or3_4
Xhold1303 _15346_/D _08461_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1325 hold1325/X _15585_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 hold1314/X _15608_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08843_ VGND VPWR VPWR VGND _15170_/D _09686_/A0 _08850_/S hold562/X sky130_fd_sc_hd__mux2_1
Xhold1336 hold1336/X _15332_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1358 hold1358/X _15429_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08774_ VGND VPWR VPWR VGND _15232_/D _09862_/A0 _08779_/S hold221/X sky130_fd_sc_hd__mux2_1
Xhold1347 _08782_/A _15226_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07725_ VGND VPWR VPWR VGND _15560_/Q _07958_/A _07725_/B sky130_fd_sc_hd__xor2_1
Xhold1369 _09731_/A _14314_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07656_ VPWR VGND VPWR VGND _07668_/B _15092_/Q _07881_/A2 _07656_/X _07338_/A sky130_fd_sc_hd__a22o_1
X_07587_ VPWR VGND VPWR VGND _09007_/B _11284_/B _09010_/B _07587_/B sky130_fd_sc_hd__or3b_2
XFILLER_41_738 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09326_ VGND VPWR VPWR VGND _14718_/D hold762/X _09327_/S fanout41/X sky130_fd_sc_hd__mux2_1
X_09257_ VGND VPWR VPWR VGND _14786_/D fanout40/X _09272_/S hold493/X sky130_fd_sc_hd__mux2_1
X_13866__983 VPWR VGND VPWR VGND _15238_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
Xclone47 VPWR VGND clone47/X clone47/A VPWR VGND sky130_fd_sc_hd__buf_6
X_08208_ VPWR VGND VGND VPWR _08208_/X _08208_/A _08208_/B sky130_fd_sc_hd__or2_1
XFILLER_5_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09188_ VGND VPWR VPWR VGND _14903_/D hold644/X _09188_/S fanout7/X sky130_fd_sc_hd__mux2_1
X_08139_ VPWR VGND VGND VPWR _08139_/X _08277_/S _10062_/C sky130_fd_sc_hd__or2_1
X_13409__526 VPWR VGND VPWR VGND _14684_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_11150_ VPWR VGND VGND VPWR _11150_/X hold263/A _11251_/B sky130_fd_sc_hd__or2_1
X_10101_ VGND VPWR VPWR VGND _10101_/X hold878/A _10516_/S hold464/A sky130_fd_sc_hd__mux2_1
X_11081_ VPWR VGND VGND VPWR _11062_/Y _11080_/X _12677_/A2 _14405_/Q _14405_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
X_10032_ VPWR VGND VPWR VGND _10031_/C hold1458/X hold1304/X _10033_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_1367 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14840_ _14840_/Q clkload28/A _14840_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14771_ hold673/A _14771_/CLK _14771_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11983_ VGND VPWR VPWR VGND _11987_/B hold601/A _11998_/S hold360/A sky130_fd_sc_hd__mux2_1
X_10934_ VGND VPWR VPWR VGND _10938_/B hold567/A _11179_/S hold559/A sky130_fd_sc_hd__mux2_1
X_10865_ VGND VPWR VPWR VGND _10865_/X _14560_/Q _10885_/S hold254/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12604_ VGND VPWR VPWR VGND _12608_/B hold629/A _12623_/S hold388/A sky130_fd_sc_hd__mux2_1
X_15323_ _15323_/Q _15323_/CLK _15323_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10796_ VGND VPWR VPWR VGND _10796_/X _10795_/X _11213_/S _10794_/X sky130_fd_sc_hd__mux2_1
X_12535_ VGND VPWR VGND VPWR _12535_/X _12662_/A1 _12531_/X _12534_/X _12662_/C1 sky130_fd_sc_hd__o211a_1
X_15254_ _15254_/Q _15254_/CLK _15254_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12466_ VGND VPWR VPWR VGND _12466_/X _14211_/Q _12479_/S hold600/A sky130_fd_sc_hd__mux2_1
X_11417_ VGND VPWR VGND VPWR _14843_/Q _11368_/A _14854_/Q _11367_/D _11361_/X _11417_/X
+ sky130_fd_sc_hd__a311o_1
X_14205_ _14205_/Q _14205_/CLK _14205_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12397_ VPWR VGND VPWR VGND _12396_/X _12722_/A1 _12395_/X _12397_/Y sky130_fd_sc_hd__a21oi_1
X_15185_ hold428/A _15185_/CLK _15185_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11348_ VGND VPWR VPWR VGND _11348_/X _14926_/Q _11355_/S hold1210/X sky130_fd_sc_hd__mux2_1
X_14136_ _14136_/Q _14136_/CLK _14136_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_79_440 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11279_ VPWR VGND VGND VPWR _11280_/B _15442_/Q _11563_/B sky130_fd_sc_hd__or2_1
XFILLER_80_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13202__319 VPWR VGND VPWR VGND _14477_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_07510_ VGND VPWR VGND VPWR _15464_/Q _15463_/Q _15462_/Q _15461_/Q _07547_/B _07507_/B
+ sky130_fd_sc_hd__o41ai_2
X_14969_ hold777/A _14969_/CLK _14969_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_35_532 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13891__1008 VPWR VGND VPWR VGND _15263_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08490_ VPWR VGND VPWR VGND _15602_/Q _15604_/Q _15605_/Q _15603_/Q _11302_/B sky130_fd_sc_hd__or4_2
X_07441_ VPWR VGND VGND VPWR _15458_/Q _08546_/A _07714_/A sky130_fd_sc_hd__nand2_1
X_13553__670 VPWR VGND VPWR VGND _14884_/CLK clkload34/A sky130_fd_sc_hd__inv_2
Xfanout19 VPWR VGND fanout19/X _08051_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_07372_ VPWR VGND VPWR VGND _08162_/A _07372_/C _07372_/A _07372_/X sky130_fd_sc_hd__or3_1
X_09111_ VGND VPWR VPWR VGND _14984_/D hold622/X _09126_/S _07976_/X sky130_fd_sc_hd__mux2_1
X_09042_ VGND VPWR VPWR VGND _15048_/D hold595/X _09051_/S fanout37/X sky130_fd_sc_hd__mux2_1
Xhold411 hold411/X hold411/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 hold400/X hold400/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 hold444/X hold444/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold422/X hold422/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 hold433/X hold433/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 hold477/X hold477/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/X hold466/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 hold455/X hold455/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ VPWR VGND VPWR VGND _09943_/Y hold1209/X _09956_/S _14130_/D _09937_/Y sky130_fd_sc_hd__a22o_1
Xhold488 hold488/X hold488/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 hold499/X hold499/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09875_ VPWR VGND VGND VPWR _09875_/A _09875_/Y _09880_/B sky130_fd_sc_hd__nand2_1
Xhold1100 hold1100/X _15289_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 hold1122/X _15307_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 hold1133/X _14310_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ VGND VPWR VPWR VGND _15187_/D fanout62/X _08847_/S hold416/X sky130_fd_sc_hd__mux2_1
Xhold1111 hold1111/X _15002_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 hold1144/X _15432_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 hold1166/X _15701_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 hold1155/X _14758_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 _14840_/D _11353_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 hold1177/X _14502_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 hold1199/X _14438_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ VGND VPWR VPWR VGND _15249_/D _08773_/S clone46/A hold1149/X sky130_fd_sc_hd__mux2_4
X_07708_ VPWR VGND VGND VPWR _15564_/Q _07710_/A _07709_/B sky130_fd_sc_hd__nand2_1
X_08688_ VPWR VGND VPWR VGND _15284_/Q _08562_/A _08688_/X _08728_/B1 _08687_/X _08688_/C1
+ sky130_fd_sc_hd__a221o_1
X_07639_ VPWR VGND VGND VPWR _07639_/A _07859_/B _07639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10650_ VPWR VGND VGND VPWR _10650_/X _10652_/S _10650_/B sky130_fd_sc_hd__or2_1
X_09309_ VGND VPWR VPWR VGND _14732_/D fanout98/X _09310_/S hold309/X sky130_fd_sc_hd__mux2_1
XFILLER_16_1013 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10581_ VPWR VGND VGND VPWR _10729_/A _10581_/B _10581_/Y sky130_fd_sc_hd__nor2_1
X_12320_ VPWR VGND VGND VPWR _12320_/X _12684_/S _12320_/B sky130_fd_sc_hd__or2_1
X_12251_ VGND VPWR VPWR VGND _12251_/X hold808/A _12578_/S hold581/A sky130_fd_sc_hd__mux2_1
X_11202_ VGND VPWR VPWR VGND _11202_/X hold557/A _11204_/S hold323/A sky130_fd_sc_hd__mux2_1
XFILLER_79_88 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12182_ VGND VPWR VGND VPWR _12182_/X hold992/A _12192_/A2 _11958_/A _12181_/X sky130_fd_sc_hd__o211a_1
X_11133_ VGND VPWR VPWR VGND _11133_/X _11130_/X _11143_/S _11129_/X sky130_fd_sc_hd__mux2_1
X_14053__1170 VPWR VGND VPWR VGND _15425_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_11064_ VGND VPWR VPWR VGND _11064_/X hold783/A _11175_/S hold708/A sky130_fd_sc_hd__mux2_1
X_10015_ VPWR VGND VGND VPWR _10017_/C _10015_/B _15621_/D sky130_fd_sc_hd__nor2_1
X_13496__613 VPWR VGND VPWR VGND _14771_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
XFILLER_0_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14823_ hold147/A clkload29/A input4/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_28_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11966_ VPWR VGND VGND VPWR _11966_/X _12164_/A _11966_/B sky130_fd_sc_hd__or2_1
X_13537__654 VPWR VGND VPWR VGND _14868_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_14754_ hold251/A _14754_/CLK _14754_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14685_ hold684/A _14685_/CLK _14685_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10917_ VGND VPWR VPWR VGND _10917_/X hold831/A _10924_/B _14916_/Q sky130_fd_sc_hd__mux2_1
X_11897_ VPWR VGND _11897_/X _11871_/X _11867_/X _12111_/C1 _12029_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_10848_ VGND VPWR VPWR VGND _10848_/X _15019_/Q _11107_/S hold757/A sky130_fd_sc_hd__mux2_1
X_10779_ VPWR VGND VGND VPWR _10779_/X hold311/A _10850_/S sky130_fd_sc_hd__or2_1
X_15306_ _15306_/Q _15306_/CLK _15306_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12938__55 VPWR VGND VPWR VGND _14181_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_12518_ VGND VPWR VGND VPWR _12518_/X _12656_/A1 _12513_/X _12517_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_15237_ hold177/A _15237_/CLK _15237_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12449_ VPWR VGND VGND VPWR _12449_/X hold156/A _12623_/S sky130_fd_sc_hd__or2_1
X_15168_ hold523/A _15168_/CLK _15168_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15099_ _15099_/Q _15099_/CLK _15099_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07990_ VPWR VGND VGND VPWR _07990_/X _07990_/A _07990_/B sky130_fd_sc_hd__or2_1
Xfanout209 VGND VPWR _12674_/A1 _12737_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_80_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09660_ VPWR VGND VPWR VGND _09660_/X _09764_/A _09660_/B sky130_fd_sc_hd__or2_2
X_14210__928 _14210_/D _14210__928/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xtt_um_femto_903 uio_out[6] tt_um_femto_903/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08611_ VPWR VGND VGND VPWR _08617_/A _09004_/B _08611_/Y sky130_fd_sc_hd__nor2_1
X_09591_ VPWR VGND VGND VPWR _09591_/Y _09764_/A _09591_/A sky130_fd_sc_hd__nor2_4
X_08542_ VPWR VGND VGND VPWR _15558_/Q _08542_/Y _09976_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_1084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08473_ VGND VPWR VGND VPWR _15340_/D hold1190/X _08483_/A2 _08472_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_1024 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07424_ VPWR VGND VGND VPWR _07424_/X _07974_/B1 _07423_/X _07419_/X _07416_/Y _07413_/Y
+ sky130_fd_sc_hd__o41a_1
X_07355_ VPWR VGND VGND VPWR _11973_/A _07355_/B _07355_/Y sky130_fd_sc_hd__nor2_1
X_13330__447 VPWR VGND VPWR VGND _14605_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_07286_ VPWR VGND VPWR VGND _07925_/A _07926_/A _07286_/B sky130_fd_sc_hd__or2_2
X_09025_ VPWR VGND VPWR VGND _09022_/B _09974_/A _15063_/D _09024_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_40_49 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold252 hold252/X hold252/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/X hold230/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13183__300 VPWR VGND VPWR VGND _14458_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
Xhold241 hold241/X hold241/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/X hold274/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/X hold296/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/X hold285/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/X hold263/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 VGND VPWR _08424_/Y _08484_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09927_ VGND VPWR VPWR VGND _14135_/D hold1206/X _09931_/B _09926_/X sky130_fd_sc_hd__mux2_1
Xfanout721 VGND VPWR _11974_/A1 _12195_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout732 VPWR VGND _12751_/A2 _12269_/B VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout743 VGND VPWR _07828_/Y _07886_/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout765 VPWR VGND _08002_/A2 _07425_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout754 VGND VPWR _07826_/X _12790_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout776 VGND VPWR _08225_/C1 _08280_/B2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13224__341 VPWR VGND VPWR VGND _14499_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
Xfanout787 VPWR VGND _09938_/A _07534_/A VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout798 VPWR VGND _08617_/A _08582_/A VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_63_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09858_ VGND VPWR VPWR VGND _14164_/D hold453/X _09865_/S fanout7/X sky130_fd_sc_hd__mux2_1
X_08809_ VGND VPWR VPWR VGND _15200_/D _09862_/A0 _08814_/S hold404/X sky130_fd_sc_hd__mux2_1
X_09789_ VGND VPWR VPWR VGND _14260_/D fanout7/X _09790_/S hold730/X sky130_fd_sc_hd__mux2_1
XANTENNA_114 _09161_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11820_ VGND VPWR VPWR VGND _11820_/X hold797/A _12372_/S hold495/A sky130_fd_sc_hd__mux2_1
XANTENNA_103 _10846_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11751_ VPWR VGND VPWR VGND _11750_/X _12473_/A _12491_/B1 _11751_/X sky130_fd_sc_hd__a21o_1
X_10702_ VGND VPWR VPWR VGND _10702_/X hold528/A _10702_/S hold270/A sky130_fd_sc_hd__mux2_1
X_14470_ _14470_/Q _14470_/CLK _14470_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11682_ VGND VPWR VPWR VGND _11682_/X hold503/A _12052_/S hold219/A sky130_fd_sc_hd__mux2_1
X_13962__1079 VPWR VGND VPWR VGND _15334_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_10633_ VGND VPWR VGND VPWR _10633_/X _15013_/Q _10633_/A2 _10632_/X _10625_/S sky130_fd_sc_hd__o211a_1
X_10564_ VGND VPWR VPWR VGND _10568_/B hold760/A _10730_/S hold654/A sky130_fd_sc_hd__mux2_1
XFILLER_10_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12303_ VGND VPWR VPWR VGND _12303_/X hold568/A _12708_/S hold261/A sky130_fd_sc_hd__mux2_1
XFILLER_6_734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10495_ VGND VPWR VGND VPWR _10495_/X _10523_/A1 _10491_/X _10494_/X _10630_/C1 sky130_fd_sc_hd__o211a_1
X_15022_ _15022_/Q _15022_/CLK _15022_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12234_ VGND VPWR VPWR VGND _12234_/X hold619/A _12578_/S hold376/A sky130_fd_sc_hd__mux2_1
X_13890__1007 VPWR VGND VPWR VGND _15262_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_12165_ VGND VPWR VGND VPWR _12165_/X _11958_/A _12161_/X _12164_/X _12184_/C1 sky130_fd_sc_hd__o211a_1
X_11116_ VPWR VGND VPWR VGND _11116_/X _11173_/A _11089_/X _11097_/X _11115_/X _11114_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_7_1044 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12096_ VGND VPWR VPWR VGND _12096_/X _14201_/Q _12097_/S _15209_/Q sky130_fd_sc_hd__mux2_1
X_11047_ VGND VPWR VPWR VGND _11047_/X hold946/A _11054_/S hold893/A sky130_fd_sc_hd__mux2_1
X_14806_ _14806_/Q _14806_/CLK _14806_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13771__888 VPWR VGND VPWR VGND _15143_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_79_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14737_ hold163/A _14737_/CLK _14737_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11949_ VGND VPWR VPWR VGND _11949_/X hold879/A _11950_/B hold189/A sky130_fd_sc_hd__mux2_1
X_14668_ hold702/A _14668_/CLK _14668_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_696 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07140_ VPWR VGND VGND VPWR _07826_/A _15574_/Q wire858/A _15572_/Q _07765_/B sky130_fd_sc_hd__nor4b_1
X_14599_ hold326/A _14599_/CLK _14599_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13665__782 VPWR VGND VPWR VGND _15005_/CLK clkload49/A sky130_fd_sc_hd__inv_2
X_13208__325 VPWR VGND VPWR VGND _14483_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_09712_ VGND VPWR VPWR VGND _14331_/D fanout31/X _09728_/S hold938/X sky130_fd_sc_hd__mux2_1
X_07973_ VPWR VGND VPWR VGND _15082_/Q _10072_/B _07973_/X _10074_/A0 _07182_/A _07972_/Y
+ sky130_fd_sc_hd__a221o_1
XFILLER_56_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09643_ VGND VPWR VPWR VGND _14427_/D hold998/X _09659_/S fanout33/X sky130_fd_sc_hd__mux2_1
X_09574_ VGND VPWR VPWR VGND _14491_/D hold1006/X _09590_/S fanout32/X sky130_fd_sc_hd__mux2_1
X_08525_ VGND VPWR VGND VPWR _15324_/D hold1216/X _08553_/A2 _08524_/Y _11398_/A sky130_fd_sc_hd__o211a_1
XFILLER_58_1422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_62_clk clkload18/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_08456_ VPWR VGND VGND VPWR _08456_/X _15348_/Q _08486_/B sky130_fd_sc_hd__or2_1
X_07407_ VPWR VGND VGND VPWR _07607_/B _07607_/C _07612_/A _07410_/C sky130_fd_sc_hd__o21a_1
X_08387_ VGND VPWR VPWR VGND _15390_/D fanout62/X _08408_/S hold810/X sky130_fd_sc_hd__mux2_1
X_07338_ VPWR VGND VPWR VGND _07653_/A _07338_/A _07338_/B sky130_fd_sc_hd__or2_2
XFILLER_13_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07269_ VPWR VGND VPWR VGND _08025_/A _08026_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09008_ VGND VPWR VGND VPWR _09008_/X _09007_/A _09016_/B1 _15100_/Q _09007_/Y sky130_fd_sc_hd__a211o_1
X_10280_ VPWR VGND VGND VPWR _10280_/X _10613_/A _10280_/B sky130_fd_sc_hd__or2_1
Xfanout551 VPWR VGND clone13/A _07557_/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout540 VPWR VGND _08711_/B1 _08662_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout573 _09411_/S _09381_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout562 VPWR VGND _09659_/S _09657_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout584 VPWR VGND _09157_/S _09160_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout595 VGND VPWR _08816_/Y _08847_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15640_ VGND VPWR VPWR VGND _15640_/Q _15640_/D _10060_/Y sky130_fd_sc_hd__dlxtn_1
X_12852_ VGND VPWR VPWR VGND _15576_/D _08176_/X _12860_/S _12878_/A sky130_fd_sc_hd__mux2_1
X_13001__118 VPWR VGND VPWR VGND _14244_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_11803_ VGND VPWR VGND VPWR _11803_/X _12588_/A1 _11799_/X _11802_/X _12748_/C1 sky130_fd_sc_hd__o211a_1
X_12783_ VPWR VGND VGND VPWR _12790_/A _12783_/Y _12783_/B sky130_fd_sc_hd__nand2_1
X_15571_ _15571_/Q clkload15/A _15571_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_53_clk _12980__97/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_42_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11734_ VGND VPWR VPWR VGND _11734_/X hold839/A _12409_/B hold638/A sky130_fd_sc_hd__mux2_1
X_14522_ hold241/A _14522_/CLK _14522_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11665_ VGND VPWR VPWR VGND _11665_/X hold927/A _11964_/S hold445/A sky130_fd_sc_hd__mux2_1
X_14453_ hold596/A _14453_/CLK _14453_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10616_ VPWR VGND VPWR VGND _10615_/X _10616_/A1 _10614_/X _10616_/Y sky130_fd_sc_hd__a21oi_1
X_13649__766 VPWR VGND VPWR VGND _14989_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_11596_ VGND VPWR VGND VPWR _11596_/X _14999_/Q _12040_/A2 _11625_/S _11595_/X sky130_fd_sc_hd__o211a_1
X_14384_ VGND VPWR VGND VPWR _14384_/Q _14384_/D clkload11/A sky130_fd_sc_hd__dfxtp_4
X_12908__25 VPWR VGND VPWR VGND _14150_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_10547_ VGND VPWR VPWR VGND _10547_/X hold637/A _10627_/S hold858/A sky130_fd_sc_hd__mux2_1
X_10478_ VGND VPWR VGND VPWR _10478_/X _10706_/C1 _10473_/X _10477_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_15005_ _15005_/Q _15005_/CLK _15005_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12217_ VGND VPWR VPWR VGND _12217_/X hold792/A _12228_/B hold466/A sky130_fd_sc_hd__mux2_1
X_12148_ VGND VPWR VGND VPWR _12148_/X _12212_/A1 _12147_/X _12144_/X _12222_/C1 sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12079_ VPWR VGND VGND VPWR _12079_/X hold155/A _12227_/S sky130_fd_sc_hd__or2_1
XFILLER_38_925 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_80_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_928 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_clk clkload38/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09290_ VGND VPWR VPWR VGND _14751_/D fanout47/X _09304_/S hold217/X sky130_fd_sc_hd__mux2_1
X_08310_ VGND VPWR VPWR VGND _15509_/D fanout77/X _08318_/S hold824/X sky130_fd_sc_hd__mux2_1
X_08241_ VGND VPWR VPWR VGND _10062_/A _08241_/X _08241_/B sky130_fd_sc_hd__xor2_1
XANTENNA_14 _09061_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_25 _14402_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_47 _08178_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_36 _12864_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XANTENNA_69 _09865_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08172_ VGND VPWR VPWR VGND _08172_/X _07331_/A _08195_/A _08232_/B _08197_/S sky130_fd_sc_hd__o31a_2
X_14032__1149 VPWR VGND VPWR VGND _15404_/CLK clkload55/A sky130_fd_sc_hd__inv_2
XANTENNA_58 fanout539/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07123_ VPWR VGND VPWR VGND _07123_/Y _07123_/A sky130_fd_sc_hd__inv_2
XFILLER_0_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14216__934 _14216_/D _14216__934/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_13442__559 VPWR VGND VPWR VGND _14717_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_13961__1078 VPWR VGND VPWR VGND _15333_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_07956_ VPWR VGND VPWR VGND clone19/X _15349_/Q clone13/X _07956_/X _15138_/Q sky130_fd_sc_hd__a22o_1
XFILLER_25_1421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07887_ VPWR VGND VPWR VGND _15627_/Q _07952_/A2 _07890_/A _07908_/B1 _15591_/Q _07886_/Y
+ sky130_fd_sc_hd__a221o_1
X_13295__412 VPWR VGND VPWR VGND _14570_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_09626_ VGND VPWR VGND VPWR _09660_/B _09694_/A _09626_/X sky130_fd_sc_hd__or2_4
X_09557_ VPWR VGND VGND VPWR _09557_/Y _09557_/A _09834_/B sky130_fd_sc_hd__nand2_2
X_08508_ VGND VPWR VPWR VGND _08508_/B _08507_/C _08508_/A _08508_/X sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_35_clk _12964__81/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_13336__453 VPWR VGND VPWR VGND _14611_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_09488_ VPWR VGND VGND VPWR _09488_/X _09488_/A _09517_/S sky130_fd_sc_hd__or2_1
XFILLER_19_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08439_ VGND VPWR VGND VPWR _15357_/D _15356_/Q _08448_/B _08438_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_51_482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11450_ VGND VPWR VPWR VGND _15067_/D _11449_/X _11480_/S hold1391/X sky130_fd_sc_hd__mux2_1
XFILLER_32_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11381_ VGND VPWR VPWR VGND _11381_/X _11380_/X _11387_/S _14848_/Q sky130_fd_sc_hd__mux2_1
X_10401_ VGND VPWR VGND VPWR _10401_/X hold835/A _10688_/A2 _10400_/X _10698_/A1 sky130_fd_sc_hd__o211a_1
X_10332_ VGND VPWR VPWR VGND _10332_/X hold398/A _11098_/S hold235/A sky130_fd_sc_hd__mux2_1
X_12002_ VGND VPWR VGND VPWR _12002_/X hold802/A _12188_/A2 _12008_/A1 _12001_/X sky130_fd_sc_hd__o211a_1
X_10263_ VGND VPWR VGND VPWR _10263_/X _15003_/Q _11003_/A2 _10262_/X _11244_/S sky130_fd_sc_hd__o211a_1
X_10194_ VGND VPWR VPWR VGND _10198_/B hold368/A _10972_/S hold635/A sky130_fd_sc_hd__mux2_1
XFILLER_78_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout370 VPWR VGND _10333_/A fanout382/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout381 VPWR VGND fanout381/X fanout382/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_4_1014 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout392 VGND VPWR _10593_/A1 _10745_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_35_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12835_ VPWR VGND VPWR VGND _12833_/X _15566_/Q _10056_/Y _15566_/D _12834_/X sky130_fd_sc_hd__a22o_1
X_15623_ _15623_/Q clkload50/A _15623_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15554_ _15554_/Q clkload32/A _15554_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_26_clk clkload43/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_76_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14505_ hold903/A _14505_/CLK _14505_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12766_ VPWR VGND VGND VPWR _12766_/X _12822_/A _12766_/B sky130_fd_sc_hd__or2_1
X_13079__196 VPWR VGND VPWR VGND _14322_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_12697_ VGND VPWR VPWR VGND _12697_/X hold980/A _12701_/S hold911/A sky130_fd_sc_hd__mux2_1
X_11717_ VGND VPWR VPWR VGND _11717_/X hold968/A _11748_/S hold731/A sky130_fd_sc_hd__mux2_1
X_15485_ _15485_/Q _15485_/CLK _15485_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11648_ VGND VPWR VPWR VGND _11648_/X _11645_/X _11948_/S _11644_/X sky130_fd_sc_hd__mux2_1
X_14436_ hold925/A _14436_/CLK _14436_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14367_ hold880/A _14367_/CLK _14367_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11579_ VGND VPWR VPWR VGND _11579_/X hold789/A _12086_/S hold165/A sky130_fd_sc_hd__mux2_1
Xhold807 hold807/X hold807/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold818 hold818/X hold818/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_862 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold829 hold829/X hold829/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ hold621/A _14298_/CLK _14298_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07810_ VPWR VGND _07849_/A _07810_/B _07810_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08790_ VGND VPWR VPWR VGND _15219_/D fanout60/X _08811_/S hold600/X sky130_fd_sc_hd__mux2_1
XFILLER_78_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13777__894 VPWR VGND VPWR VGND _15149_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_07741_ VPWR VGND _07741_/X _07742_/B _15554_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_42_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07672_ VPWR VGND VPWR VGND _15632_/Q _07952_/A2 _07673_/B _07908_/B1 _15596_/Q _07671_/Y
+ sky130_fd_sc_hd__a221o_1
X_13023__140 VPWR VGND VPWR VGND _14266_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_0_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09411_ VGND VPWR VPWR VGND _14638_/D hold635/X _09411_/S _09864_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_20_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_17_clk _12891__8/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09342_ VGND VPWR VPWR VGND _14702_/D hold468/X _09342_/S _09690_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_34_994 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_482 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09273_ VGND VPWR VPWR VGND _14770_/D _09865_/A0 _09275_/S hold666/X sky130_fd_sc_hd__mux2_1
X_08224_ VPWR VGND VPWR VGND _08223_/Y _08201_/C _08240_/A _08224_/X sky130_fd_sc_hd__a21o_1
X_08155_ VPWR VGND VGND VPWR _08155_/X _08155_/A _08155_/B sky130_fd_sc_hd__or2_1
X_07106_ VPWR VGND VPWR VGND _07106_/Y _14858_/Q sky130_fd_sc_hd__inv_2
X_08086_ VPWR VGND VPWR VGND _08293_/A3 _07190_/B _08278_/B _08086_/X _07188_/X sky130_fd_sc_hd__a22o_1
X_12899__16 VPWR VGND VPWR VGND _14141_/CLK clkload29/A sky130_fd_sc_hd__inv_2
XFILLER_62_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08988_ VGND VPWR VGND VPWR _15108_/D hold1056/X _09015_/A2 _08987_/X _11337_/C1
+ sky130_fd_sc_hd__o211a_1
X_07939_ VGND VPWR _07939_/B _07939_/Y _07939_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_10950_ VGND VPWR VPWR VGND _10951_/B _10949_/Y _11246_/S _10941_/Y sky130_fd_sc_hd__mux2_1
XFILLER_17_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_71_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10881_ VGND VPWR VPWR VGND _10881_/X hold769/A _10885_/S hold475/A sky130_fd_sc_hd__mux2_1
X_09609_ VGND VPWR VPWR VGND _14459_/D fanout31/X _09625_/S hold694/X sky130_fd_sc_hd__mux2_1
XFILLER_73_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12620_ VGND VPWR VPWR VGND _12621_/B _12619_/Y _12731_/S _12611_/Y sky130_fd_sc_hd__mux2_1
X_13570__687 VPWR VGND VPWR VGND _14901_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_12551_ VGND VPWR VGND VPWR _12551_/X _12550_/X _12549_/X _12670_/A1 _12670_/C1 sky130_fd_sc_hd__a211o_1
X_11502_ VGND VPWR VPWR VGND _11502_/X _15086_/Q _11535_/C _15084_/Q sky130_fd_sc_hd__mux2_1
X_15270_ hold977/A _15270_/CLK _15270_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12482_ VGND VPWR VPWR VGND _12482_/X hold810/A _12716_/S hold204/A sky130_fd_sc_hd__mux2_1
X_11433_ VGND VPWR VGND VPWR _14931_/D _14932_/Q _11439_/A2 _11432_/X _09977_/A sky130_fd_sc_hd__o211a_1
X_14221_ hold257/A _14221_/CLK _14221_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14152_ hold212/A _14152_/CLK _14152_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11364_ VGND VPWR VPWR VGND _11364_/X _14843_/Q _11392_/B _14811_/Q sky130_fd_sc_hd__mux2_1
X_10315_ VGND VPWR VPWR VGND _10315_/X _10314_/X _10315_/S _10313_/X sky130_fd_sc_hd__mux2_1
X_11295_ VGND VPWR VPWR VGND _11296_/B _14816_/Q _11299_/S _14384_/Q sky130_fd_sc_hd__mux2_1
XFILLER_3_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13464__581 VPWR VGND VPWR VGND _14739_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_10246_ VPWR VGND VPWR VGND _10245_/X _10930_/C1 _10244_/X _10246_/Y sky130_fd_sc_hd__a21oi_1
X_10177_ VGND VPWR VPWR VGND _10177_/X hold948/A _10472_/S hold649/A sky130_fd_sc_hd__mux2_1
X_14985_ hold685/A _14985_/CLK _14985_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14031__1148 VPWR VGND VPWR VGND _15403_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_13007__124 VPWR VGND VPWR VGND _14250_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_13811__928 VPWR VGND VPWR VGND _15183_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_15606_ hold807/A clkload27/A _15606_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12818_ VPWR VGND VPWR VGND _07918_/Y _12790_/A _09975_/A _12818_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12749_ VPWR VGND _12749_/X _12748_/X _12744_/X _12583_/S _12740_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15537_ hold204/A _15537_/CLK _15537_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15468_ _15468_/Q clkload41/A _15468_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_13960__1077 VPWR VGND VPWR VGND _15332_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_14419_ hold933/A _14419_/CLK _14419_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_485 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15399_ hold345/A _15399_/CLK _15399_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold615 hold615/X hold615/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 hold604/X hold604/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13705__822 VPWR VGND VPWR VGND _15045_/CLK clkload10/A sky130_fd_sc_hd__inv_2
Xhold626 hold626/X hold626/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ VPWR VGND VGND VPWR hold148/X _08502_/B _08529_/A _14765_/D sky130_fd_sc_hd__o21a_1
Xhold659 hold659/X hold659/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clkload10/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold637 hold637/X hold637/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 hold648/X hold648/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08911_ VGND VPWR VGND VPWR _15137_/D hold1279/X _08919_/A2 _08910_/X _08919_/C1
+ sky130_fd_sc_hd__o211a_1
X_09891_ VGND VPWR VPWR VGND _09892_/C _07123_/Y _09891_/S _09970_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_839 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08842_ VGND VPWR VPWR VGND _15171_/D _09685_/A0 _08842_/S hold399/X sky130_fd_sc_hd__mux2_1
Xhold1304 hold1304/X _15629_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1315 _09984_/B _09983_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 _09916_/A _14138_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1337 _15333_/D _08487_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1359 hold1359/X _14134_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08773_ VGND VPWR VPWR VGND _15233_/D _09827_/A1 _08773_/S hold279/X sky130_fd_sc_hd__mux2_1
Xhold1348 _10007_/A _15618_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07724_ VPWR VGND _07800_/A _07725_/B _15560_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07655_ _07655_/X _07857_/A _07649_/Y _07650_/X _07654_/Y _10071_/A VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__o311a_1
X_07586_ VPWR VGND VGND VPWR _08174_/A _09007_/B _07586_/C _11302_/A sky130_fd_sc_hd__nor3_2
X_09325_ VGND VPWR VPWR VGND _14719_/D hold652/X _09342_/S fanout44/X sky130_fd_sc_hd__mux2_1
XFILLER_22_953 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09256_ VGND VPWR VPWR VGND _14787_/D clone44/A _09272_/S hold438/X sky130_fd_sc_hd__mux2_1
X_08207_ VPWR VGND VGND VPWR _15548_/Q _08220_/B _08208_/B sky130_fd_sc_hd__nor2_1
X_09187_ VGND VPWR VPWR VGND _14904_/D hold356/X _09197_/S fanout8/X sky130_fd_sc_hd__mux2_1
XFILLER_5_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08138_ VPWR VGND VGND VPWR _08138_/A _08138_/B _10062_/C sky130_fd_sc_hd__nor2_1
X_13448__565 VPWR VGND VPWR VGND _14723_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XFILLER_49_1048 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08069_ _08070_/D _08065_/X _08066_/Y _08068_/X _08294_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_66_1351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11080_ VPWR VGND VPWR VGND _11079_/X _11247_/A _12713_/B1 _11080_/X sky130_fd_sc_hd__a21o_1
X_10100_ VPWR VGND VGND VPWR _10618_/A _10100_/B _10100_/Y sky130_fd_sc_hd__nor2_1
X_10031_ VGND VPWR _10035_/B _15629_/Q _15628_/Q _10031_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_1_857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14770_ hold666/A _14770_/CLK _14770_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11982_ VPWR VGND VPWR VGND _11981_/X _12008_/C1 _11980_/X _11982_/Y sky130_fd_sc_hd__a21oi_1
X_10933_ VPWR VGND VGND VPWR _10914_/Y _10932_/X _12751_/A2 _14401_/Q _14401_/D _12751_/C1
+ sky130_fd_sc_hd__o221a_1
X_10864_ VGND VPWR VGND VPWR _10864_/X hold973/A _12866_/A1 _10863_/X _10890_/A sky130_fd_sc_hd__o211a_1
X_12603_ VPWR VGND VGND VPWR _12584_/Y _12602_/X _12269_/B _15472_/Q _15472_/D _11341_/A
+ sky130_fd_sc_hd__o221a_1
X_10795_ VGND VPWR VPWR VGND _10795_/X hold378/A _10795_/S hold620/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15322_ _15322_/Q _15322_/CLK _15322_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12534_ VPWR VGND VGND VPWR _12534_/X _12665_/S _12534_/B sky130_fd_sc_hd__or2_1
XFILLER_33_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15253_ hold893/A _15253_/CLK _15253_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12465_ VGND VPWR VPWR VGND _12465_/X hold507/A _12479_/S hold293/A sky130_fd_sc_hd__mux2_1
X_11416_ VPWR VGND _14859_/D _11415_/X _11368_/A _08541_/A _11396_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15184_ _15184_/Q _15184_/CLK _15184_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12396_ VGND VPWR VPWR VGND _12396_/X _12393_/X _12396_/S _12392_/X sky130_fd_sc_hd__mux2_1
X_14204_ _14204_/Q _14204_/CLK _14204_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11347_ VGND VPWR _14834_/D _11347_/B _11347_/A _11347_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14135_ _14135_/Q _14135_/CLK _14135_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11278_ VPWR VGND VGND VPWR _11563_/B _15441_/Q _11561_/B sky130_fd_sc_hd__or2_1
XFILLER_45_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10229_ VPWR VGND VPWR VGND _10228_/X _11210_/A _12491_/B1 _10229_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13241__358 VPWR VGND VPWR VGND _14516_/CLK clkload17/A sky130_fd_sc_hd__inv_2
XFILLER_47_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14968_ hold549/A _14968_/CLK _14968_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14899_ hold362/A _14899_/CLK _14899_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07440_ VPWR VGND VGND VPWR _08554_/A _08548_/B _07440_/B sky130_fd_sc_hd__or2_1
XFILLER_50_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13094__211 VPWR VGND VPWR VGND _14337_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07371_ VPWR VGND VGND VPWR _07371_/X _07371_/A _07371_/B sky130_fd_sc_hd__or2_1
X_09110_ VGND VPWR VPWR VGND _14985_/D hold685/X _09122_/S fanout38/X sky130_fd_sc_hd__mux2_1
X_09041_ VGND VPWR VPWR VGND _15049_/D hold432/X _09053_/S fanout38/X sky130_fd_sc_hd__mux2_1
X_13135__252 VPWR VGND VPWR VGND _14378_/CLK clkload39/A sky130_fd_sc_hd__inv_2
Xhold401 hold401/X hold401/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 hold445/X hold445/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 hold412/X hold412/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 hold423/X hold423/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 hold434/X hold434/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 hold478/X hold478/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 hold467/X hold467/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 hold456/X hold456/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ VPWR VGND VGND VPWR _09947_/C _09943_/Y _09943_/B sky130_fd_sc_hd__nand2_1
Xhold489 hold489/X hold489/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09874_ VPWR VGND VGND VPWR _09878_/B _14151_/Q _09880_/B sky130_fd_sc_hd__or2_1
Xhold1123 hold1123/X _14182_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 hold1112/X _15000_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ VGND VPWR VPWR VGND _15188_/D fanout64/X _08846_/S hold775/X sky130_fd_sc_hd__mux2_1
Xhold1101 hold1101/X _15004_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 hold1145/X _14144_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _14861_/D _11420_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 hold1156/X _15425_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 hold1134/X _15491_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1189 hold1189/X _14789_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 hold1178/X _15387_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13833__950 VPWR VGND VPWR VGND _15205_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_08756_ VGND VPWR VPWR VGND _08773_/S fanout57/X hold1141/X _15250_/D sky130_fd_sc_hd__mux2_2
X_12999__116 VPWR VGND VPWR VGND _14242_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_07707_ VGND VPWR VPWR VGND _07709_/B _15591_/Q _07807_/S _07519_/B sky130_fd_sc_hd__mux2_1
X_08687_ VGND VPWR VPWR VGND _08687_/X _14396_/Q _08687_/S _14380_/Q sky130_fd_sc_hd__mux2_1
XFILLER_57_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07638_ VGND VPWR VGND VPWR _07638_/X _07966_/A _07637_/Y _07635_/X _10071_/A sky130_fd_sc_hd__o211a_1
X_07569_ VGND VPWR VGND VPWR _07567_/Y _08034_/B1 _07569_/X _15152_/Q sky130_fd_sc_hd__a21bo_4
XFILLER_53_385 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09308_ VGND VPWR VPWR VGND _14733_/D _09865_/A0 _09310_/S hold297/X sky130_fd_sc_hd__mux2_1
X_10580_ VGND VPWR VPWR VGND _10581_/B _10579_/Y _10728_/S _10571_/Y sky130_fd_sc_hd__mux2_1
X_09239_ VPWR VGND VGND VPWR hold280/X _09239_/B _14805_/D sky130_fd_sc_hd__nor2_1
X_12250_ VGND VPWR VPWR VGND _12250_/X hold868/A _12578_/S hold452/A sky130_fd_sc_hd__mux2_1
X_14030__1147 VPWR VGND VPWR VGND _15402_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_11201_ VGND VPWR VPWR VGND _11205_/B hold489/A _11204_/S hold377/A sky130_fd_sc_hd__mux2_1
X_12181_ VPWR VGND VGND VPWR _12181_/X hold337/A _12183_/S sky130_fd_sc_hd__or2_1
X_13682__799 VPWR VGND VPWR VGND _15022_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11132_ VGND VPWR VGND VPWR _11132_/X _11189_/A1 _11128_/X _11131_/X _11254_/C1 sky130_fd_sc_hd__o211a_1
Xhold990 hold990/X hold990/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ VGND VPWR VPWR VGND _11063_/X _14437_/Q _11175_/S hold436/A sky130_fd_sc_hd__mux2_1
X_10014_ VPWR VGND VGND VPWR _10014_/A _10014_/B _10015_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14822_ _14822_/Q clkload29/A hold147/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13576__693 VPWR VGND VPWR VGND _14907_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_11965_ VGND VPWR VPWR VGND _11965_/X hold718/A _11965_/S hold248/A sky130_fd_sc_hd__mux2_1
X_14753_ _14753_/Q _14753_/CLK _14753_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_17_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_555 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Right_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_60_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14684_ hold722/A _14684_/CLK _14684_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10916_ VGND VPWR VGND VPWR _10916_/X hold966/A _11003_/A2 _10915_/X _11244_/S sky130_fd_sc_hd__o211a_1
X_11896_ VGND VPWR VPWR VGND _11896_/X _11895_/X _12139_/S _11887_/X sky130_fd_sc_hd__mux2_1
X_10847_ VGND VPWR VPWR VGND _10851_/B hold501/A _11107_/S hold518/A sky130_fd_sc_hd__mux2_1
XFILLER_60_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13119__236 VPWR VGND VPWR VGND _14362_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_10778_ VGND VPWR VGND VPWR _10778_/X _10775_/X _10777_/X _11112_/A _11263_/C1 sky130_fd_sc_hd__a211o_1
X_15305_ _15305_/Q _15305_/CLK _15305_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12517_ VGND VPWR VGND VPWR _12517_/X _12516_/X _12515_/X _12665_/S _12662_/C1 sky130_fd_sc_hd__a211o_1
X_15236_ hold496/A _15236_/CLK _15236_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12448_ VGND VPWR VGND VPWR _12448_/X _12445_/X _12447_/X _12737_/B1 _12740_/A1 sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_75_Right_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12379_ VPWR VGND VGND VPWR _12360_/X _12377_/X _07913_/Y _12378_/X _12379_/X sky130_fd_sc_hd__o22a_1
X_15167_ hold609/A _15167_/CLK _15167_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15098_ _15098_/Q _15098_/CLK _15098_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_femto_904 uio_out[7] tt_um_femto_904/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08610_ VGND VPWR VPWR VGND _09004_/B _15548_/Q _07552_/B1 _10060_/C _08609_/X sky130_fd_sc_hd__o2bb2a_1
X_13817__934 VPWR VGND VPWR VGND _15189_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_28_809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09590_ VGND VPWR VPWR VGND _14475_/D hold897/X _09590_/S fanout95/X sky130_fd_sc_hd__mux2_1
X_08541_ VPWR VGND _15316_/D _08541_/B _08541_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08472_ VPWR VGND VGND VPWR _08472_/X _15340_/Q _08482_/B sky130_fd_sc_hd__or2_1
XFILLER_51_823 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07423_ VGND VPWR VPWR VGND _07423_/X _10074_/A0 _07145_/X _15476_/Q _10072_/B _15096_/Q
+ sky130_fd_sc_hd__a32o_1
XFILLER_1_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07354_ _07354_/X _07189_/B _15456_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_07285_ VPWR VGND VGND VPWR _15463_/Q _07285_/B _07946_/A sky130_fd_sc_hd__nor2_1
X_09024_ VPWR VGND VGND VPWR _09024_/A _09024_/Y _09024_/B sky130_fd_sc_hd__nand2_1
Xhold220 hold220/X hold220/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/X hold231/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/X hold242/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/X hold253/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 VGND VPWR _12870_/S _14802_/D VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold286 hold286/X hold286/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/X hold264/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/X hold275/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout733 VGND VPWR _12380_/B _12269_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09926_ VPWR VGND VPWR VGND _09925_/Y _09912_/A _08492_/X _09926_/X sky130_fd_sc_hd__a21o_1
Xhold297 hold297/X hold297/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout722 VGND VPWR _11974_/A1 _11973_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout711 VGND VPWR _08684_/S _08195_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout744 VPWR VGND _08194_/B _08233_/B VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout755 VGND VPWR _07703_/X _08147_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout766 VPWR VGND _11440_/B _08293_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
X_13263__380 VPWR VGND VPWR VGND _14538_/CLK clkload49/A sky130_fd_sc_hd__inv_2
Xfanout788 VPWR VGND _09873_/A _09890_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout799 VPWR VGND VPWR VGND _08582_/A fanout802/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09857_ VGND VPWR VPWR VGND _14165_/D hold545/X _09867_/S fanout9/X sky130_fd_sc_hd__mux2_1
Xfanout777 VGND VPWR _08225_/C1 _10071_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_08808_ VGND VPWR VPWR VGND _15201_/D _09653_/A0 _08808_/S hold243/X sky130_fd_sc_hd__mux2_1
XFILLER_58_477 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09788_ VGND VPWR VPWR VGND _14261_/D fanout9/X _09798_/S hold901/X sky130_fd_sc_hd__mux2_1
X_08739_ VGND VPWR _14764_/D _08529_/A _15261_/D _08737_/X VPWR VGND sky130_fd_sc_hd__o21ai_1
XANTENNA_115 _09864_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_104 fanout424/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11750_ VPWR VGND _11750_/X _11749_/X _11745_/X _12472_/S _11741_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10701_ VGND VPWR VPWR VGND _10705_/B hold909/A _10702_/S hold291/A sky130_fd_sc_hd__mux2_1
X_11681_ VGND VPWR VPWR VGND _11681_/X hold476/A _12052_/S hold484/A sky130_fd_sc_hd__mux2_1
X_13610__727 VPWR VGND VPWR VGND _14950_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_10632_ VPWR VGND VGND VPWR _10632_/X hold331/A _10632_/B sky130_fd_sc_hd__or2_1
X_10563_ VGND VPWR VGND VPWR _14391_/D _12121_/B1 _10561_/X _10562_/X _11294_/A sky130_fd_sc_hd__o211a_1
X_12302_ VGND VPWR VGND VPWR _12302_/X hold881/A _12746_/A2 _11810_/S _12301_/X sky130_fd_sc_hd__o211a_1
X_10494_ VPWR VGND VGND VPWR _10494_/X _10510_/S _10494_/B sky130_fd_sc_hd__or2_1
XFILLER_6_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15021_ _15021_/Q _15021_/CLK _15021_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12233_ VPWR VGND VGND VPWR _12214_/Y _12232_/X _10562_/B _15462_/Q _15462_/D _12233_/C1
+ sky130_fd_sc_hd__o221a_1
X_12164_ VPWR VGND VGND VPWR _12164_/X _12164_/A _12164_/B sky130_fd_sc_hd__or2_1
XFILLER_30_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13504__621 VPWR VGND VPWR VGND _14779_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_11115_ VPWR VGND _11115_/X _11105_/X _11101_/X _11218_/C1 _07690_/Y VGND VPWR sky130_fd_sc_hd__a31o_1
X_12095_ VGND VPWR VPWR VGND _12095_/X _14265_/Q _12097_/S hold170/A sky130_fd_sc_hd__mux2_1
X_11046_ VGND VPWR VPWR VGND _11046_/X _14501_/Q _11054_/S hold470/A sky130_fd_sc_hd__mux2_1
XFILLER_37_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14805_ hold280/A _14805_/CLK _14805_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14736_ hold390/A _14736_/CLK _14736_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11948_ VGND VPWR VPWR VGND _11948_/X _11947_/X _11948_/S _11946_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_75_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_653 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11879_ VGND VPWR VGND VPWR _11879_/X _12184_/C1 _11874_/X _11878_/X _12176_/S sky130_fd_sc_hd__o211a_1
X_14667_ hold464/A _14667_/CLK _14667_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14598_ _14598_/Q _14598_/CLK _14598_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15219_ hold600/A _15219_/CLK _15219_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13247__364 VPWR VGND VPWR VGND _14522_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_07972_ VPWR VGND VGND VPWR _07972_/A _07972_/B _07972_/Y sky130_fd_sc_hd__nor2_1
X_09711_ VGND VPWR VPWR VGND _14332_/D _07976_/X _09721_/S hold682/X sky130_fd_sc_hd__mux2_1
XFILLER_56_915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09642_ VGND VPWR VPWR VGND _14428_/D hold798/X _09657_/S fanout37/X sky130_fd_sc_hd__mux2_1
X_09573_ VGND VPWR VPWR VGND _14492_/D hold974/X _09588_/S fanout35/X sky130_fd_sc_hd__mux2_1
X_08524_ VGND VPWR _08523_/X _08553_/A2 _08524_/Y _08728_/B1 VPWR VGND sky130_fd_sc_hd__o21ai_1
X_08455_ VGND VPWR VGND VPWR _15349_/D _15348_/Q _08458_/B _08454_/X _11308_/C1 sky130_fd_sc_hd__o211a_1
X_07406_ VGND VPWR VPWR VGND _07607_/C _07343_/X _07639_/A _07625_/A _07403_/X _07665_/B
+ sky130_fd_sc_hd__o2111a_1
X_08386_ VGND VPWR VPWR VGND _15391_/D fanout64/X _08405_/S hold627/X sky130_fd_sc_hd__mux2_1
X_07337_ VPWR VGND VPWR VGND _07621_/B _07625_/A _07335_/X _07607_/B sky130_fd_sc_hd__a21o_1
XFILLER_17_1153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07268_ VPWR VGND VPWR VGND _08026_/A _07268_/A _08028_/A sky130_fd_sc_hd__or2_2
X_09007_ VPWR VGND VGND VPWR _09007_/A _09007_/B _09007_/Y sky130_fd_sc_hd__nor2_1
X_07199_ VPWR VGND VGND VPWR _07244_/A _15454_/Q _07376_/B sky130_fd_sc_hd__or2_1
Xfanout530 VGND VPWR _12594_/B _12339_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout541 VPWR VGND VPWR VGND _08662_/B1 _08522_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09909_ VPWR VGND VGND VPWR _09909_/B _09931_/B _09909_/A sky130_fd_sc_hd__nand2_4
Xfanout574 VPWR VGND _09379_/S _09377_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout552 VPWR VGND _08253_/A2 rebuffer1/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout563 VPWR VGND _09657_/S _09626_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout585 _09160_/S _09129_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_46_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout596 _08814_/S _08806_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12851_ VGND VPWR VPWR VGND _15575_/D _08193_/X _12860_/S _07328_/B sky130_fd_sc_hd__mux2_1
X_11802_ VPWR VGND VGND VPWR _11802_/X _12591_/S _11802_/B sky130_fd_sc_hd__or2_1
X_13040__157 VPWR VGND VPWR VGND _14283_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_12782_ VGND VPWR VGND VPWR _12782_/X _12788_/S _12781_/Y _08099_/Y _12790_/A sky130_fd_sc_hd__a211o_1
X_15570_ _15570_/Q clkload15/A _15570_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14521_ hold202/A _14521_/CLK _14521_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11733_ VPWR VGND VGND VPWR _12473_/A _11733_/B _11733_/Y sky130_fd_sc_hd__nor2_1
X_11664_ VGND VPWR VGND VPWR _11664_/X hold948/A _12192_/A2 _11968_/S _11663_/X sky130_fd_sc_hd__o211a_1
X_14452_ hold538/A _14452_/CLK _14452_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10615_ VGND VPWR VPWR VGND _10615_/X _10612_/X _10615_/S _10611_/X sky130_fd_sc_hd__mux2_1
X_11595_ VPWR VGND VGND VPWR _11595_/X hold532/A _11756_/S sky130_fd_sc_hd__or2_1
X_14383_ VGND VPWR VGND VPWR _14383_/Q _14383_/D clkload35/A sky130_fd_sc_hd__dfxtp_4
X_10546_ VPWR VGND VPWR VGND _10543_/X _10634_/A1 _10545_/X _10546_/X sky130_fd_sc_hd__a21o_1
X_10477_ VGND VPWR VGND VPWR _10477_/X _10476_/X _10475_/X _10467_/S _10704_/C1 sky130_fd_sc_hd__a211o_1
X_12216_ VGND VPWR VGND VPWR _12216_/X _14879_/Q _12229_/A2 _12221_/S _12215_/X sky130_fd_sc_hd__o211a_1
X_15004_ _15004_/Q _15004_/CLK _15004_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12147_ VGND VPWR VPWR VGND _12147_/X _12146_/X _12147_/S _12145_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12078_ VGND VPWR VGND VPWR _12078_/X _12075_/X _12077_/X _12230_/A1 _12230_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_65_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11029_ VGND VPWR VGND VPWR _11029_/X _11028_/X _11027_/X _11178_/C1 _11180_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_80_737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15699_ VGND VPWR hold150/A uo_out[4] VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_14719_ hold652/A _14719_/CLK _14719_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08240_ VPWR VGND VGND VPWR _08240_/A _08240_/Y _08240_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_494 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08171_ VGND VPWR VPWR VGND _15520_/D _09686_/A0 _08300_/S hold447/X sky130_fd_sc_hd__mux2_1
XANTENNA_48 _08178_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_26 _14402_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_37 _12864_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_15 _09095_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07122_ VPWR VGND VPWR VGND _09893_/A _15480_/Q sky130_fd_sc_hd__inv_2
XFILLER_53_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_59 fanout539/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_13481__598 VPWR VGND VPWR VGND _14756_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_07955_ VGND VPWR VGND VPWR _15349_/Q _07567_/B _15138_/Q _07955_/Y clone19/X sky130_fd_sc_hd__a22oi_4
XFILLER_25_1433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07886_ VPWR VGND VGND VPWR _07886_/A _07886_/B _07886_/Y sky130_fd_sc_hd__nor2_1
X_09625_ VGND VPWR VPWR VGND _14443_/D fanout97/X _09625_/S hold789/X sky130_fd_sc_hd__mux2_1
X_09556_ VPWR VGND VGND VPWR _15581_/Q _15580_/Q _09556_/C _15639_/Q _09834_/B sky130_fd_sc_hd__and4b_2
XFILLER_3_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08507_ VGND VPWR VGND VPWR _08507_/X _08507_/C _09909_/A _08508_/A sky130_fd_sc_hd__and3b_2
X_09487_ VPWR VGND VPWR VGND _09487_/Y _09517_/S sky130_fd_sc_hd__inv_2
X_13375__492 VPWR VGND VPWR VGND _14650_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_08438_ VPWR VGND VGND VPWR _08438_/X _15357_/Q _08488_/B sky130_fd_sc_hd__or2_1
X_08369_ VGND VPWR VPWR VGND _15404_/D hold315/X _08372_/S _09653_/A0 sky130_fd_sc_hd__mux2_1
X_11380_ VGND VPWR VPWR VGND _11380_/X _14847_/Q _11392_/B _14815_/Q sky130_fd_sc_hd__mux2_1
X_10400_ VPWR VGND VGND VPWR _10400_/X hold344/A _10696_/S sky130_fd_sc_hd__or2_1
X_10331_ VGND VPWR VPWR VGND _10335_/B hold782/A _11109_/S hold286/A sky130_fd_sc_hd__mux2_1
X_13722__839 VPWR VGND VPWR VGND _15062_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_10262_ VPWR VGND VGND VPWR _10262_/X hold327/A _11240_/S sky130_fd_sc_hd__or2_1
XFILLER_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12001_ VPWR VGND VGND VPWR _12001_/X hold216/A _12006_/B sky130_fd_sc_hd__or2_1
X_13929__1046 VPWR VGND VPWR VGND _15301_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_10193_ VGND VPWR VGND VPWR _14381_/D _12195_/B1 _10191_/X _10192_/X _11420_/S sky130_fd_sc_hd__o211a_1
Xfanout382 VPWR VGND fanout382/X _07873_/X VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_46_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout393 VPWR VGND _10593_/A1 fanout405/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout360 VGND VPWR _10662_/S _10652_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout371 VGND VPWR fanout381/X _11143_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13616__733 VPWR VGND VPWR VGND _14956_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_12834_ VPWR VGND VGND VPWR _12820_/B _07810_/B _12831_/A _07815_/X _12834_/X _12834_/C1
+ sky130_fd_sc_hd__o221a_1
X_15622_ _15622_/Q clkload44/A _15622_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_28_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_76_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15553_ _15553_/Q clkload31/A _15553_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12765_ VPWR VGND VGND VPWR _12822_/A _12765_/Y _12765_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11716_ VGND VPWR VPWR VGND _11720_/B hold746/A _11748_/S hold429/A sky130_fd_sc_hd__mux2_1
X_14504_ _14504_/Q _14504_/CLK _14504_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12696_ VGND VPWR VPWR VGND _12696_/X hold934/A _12701_/S hold709/A sky130_fd_sc_hd__mux2_1
X_14198__916 _14198_/D _14198__916/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_15484_ hold997/A _15484_/CLK _15484_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11647_ VGND VPWR VGND VPWR _11647_/X _11968_/S _11643_/X _11646_/X _12184_/C1 sky130_fd_sc_hd__o211a_1
X_14435_ hold939/A _14435_/CLK _14435_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14366_ hold852/A _14366_/CLK _14366_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11578_ VGND VPWR VPWR VGND _11578_/X _14187_/Q _12086_/S hold224/A sky130_fd_sc_hd__mux2_1
Xhold819 hold819/X hold819/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold808 hold808/X hold808/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ VGND VPWR VPWR VGND _10529_/X _10528_/X _10625_/S _10527_/X sky130_fd_sc_hd__mux2_1
X_14297_ hold170/A _14297_/CLK _14297_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07740_ VPWR VGND VPWR VGND _07826_/D _15590_/Q _07765_/B _07742_/B _15577_/Q sky130_fd_sc_hd__a22o_1
XFILLER_42_1087 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07671_ VPWR VGND VPWR VGND _07670_/X _07667_/X _10059_/A _07671_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13359__476 VPWR VGND VPWR VGND _14634_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_0_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09410_ VGND VPWR VPWR VGND _14639_/D hold429/X _09411_/S _09863_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_0_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09341_ VGND VPWR VPWR VGND _14703_/D hold675/X _09342_/S _09689_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_80_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_61_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09272_ VGND VPWR VPWR VGND _14771_/D _09864_/A0 _09272_/S hold673/X sky130_fd_sc_hd__mux2_1
X_08223_ VPWR VGND VGND VPWR _08223_/A _08223_/Y _08223_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12886__3 VPWR VGND VPWR VGND _14128_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08154_ VPWR VGND VPWR VGND _08208_/A _15549_/Q _15550_/Q _08155_/B sky130_fd_sc_hd__a21oi_1
XFILLER_14_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07105_ VPWR VGND VPWR VGND _09906_/A _08983_/A sky130_fd_sc_hd__inv_2
X_14810__938 _14810_/D _14810__938/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08085_ VGND VPWR VGND VPWR _08085_/X _08080_/Y _08084_/Y _08277_/S _07333_/Y sky130_fd_sc_hd__a211o_1
XFILLER_62_1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08987_ VGND VPWR VGND VPWR _08987_/X _09007_/A _09016_/B1 hold920/A _08986_/Y sky130_fd_sc_hd__a211o_1
X_13303__420 VPWR VGND VPWR VGND _14578_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_07938_ VPWR VGND VGND VPWR _07938_/A _07939_/B _07938_/B sky130_fd_sc_hd__nand2_1
X_07869_ VPWR VGND VGND VPWR _07993_/A _07869_/B _07870_/D sky130_fd_sc_hd__nor2_1
XFILLER_71_534 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10880_ VGND VPWR VPWR VGND _10880_/X _14956_/Q _10885_/S _14915_/Q sky130_fd_sc_hd__mux2_1
X_09608_ VGND VPWR VPWR VGND _14460_/D fanout35/X _09617_/S hold617/X sky130_fd_sc_hd__mux2_1
XFILLER_71_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09539_ VGND VPWR VPWR VGND _14523_/D fanout33/X _09555_/S hold291/X sky130_fd_sc_hd__mux2_1
XFILLER_52_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_40_954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12550_ VGND VPWR VPWR VGND _12550_/X hold738/A _12701_/S hold764/A sky130_fd_sc_hd__mux2_1
X_11501_ VGND VPWR VPWR VGND _15084_/D _11500_/X _11538_/S hold1395/X sky130_fd_sc_hd__mux2_1
XFILLER_11_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12481_ VGND VPWR VGND VPWR _12481_/X _12722_/A1 _12476_/X _12480_/X _12864_/A1 sky130_fd_sc_hd__o211a_1
X_11432_ VGND VPWR VGND VPWR _11432_/X _14931_/Q _11303_/A _11439_/A2 sky130_fd_sc_hd__a21bo_1
X_13152__269 VPWR VGND VPWR VGND _14427_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_14220_ hold548/A _14220_/CLK _14220_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14151_ _14151_/Q _14151_/CLK _14151_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11363_ VPWR VGND VGND VPWR _14859_/Q _14821_/Q _11406_/C sky130_fd_sc_hd__nand2b_1
XFILLER_4_844 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10314_ VGND VPWR VPWR VGND _10314_/X hold862/A _11098_/S hold163/A sky130_fd_sc_hd__mux2_1
X_11294_ VPWR VGND _14815_/D _11294_/B _11294_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_10245_ VGND VPWR VPWR VGND _10245_/X _10242_/X _10911_/S _10241_/X sky130_fd_sc_hd__mux2_1
X_10176_ VPWR VGND VPWR VGND _10173_/X _10698_/A1 _10175_/X _10176_/X sky130_fd_sc_hd__a21o_1
Xfanout190 VGND VPWR _12328_/S _11810_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13046__163 VPWR VGND VPWR VGND _14289_/CLK clkload48/A sky130_fd_sc_hd__inv_2
X_14984_ hold622/A _14984_/CLK _14984_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13850__967 VPWR VGND VPWR VGND _15222_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_12817_ VPWR VGND VGND VPWR _12817_/A _12817_/B _12817_/Y sky130_fd_sc_hd__nor2_1
X_15605_ _15605_/Q clkload19/A _15605_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12748_ VGND VPWR VGND VPWR _12748_/X _12747_/X _12746_/X _12748_/A1 _12748_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_31_932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15536_ hold162/A _15536_/CLK _15536_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12679_ VGND VPWR VPWR VGND _12679_/X hold903/A _12689_/S hold594/A sky130_fd_sc_hd__mux2_1
XFILLER_33_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15467_ _15467_/Q clkload34/A _15467_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14418_ hold919/A _14418_/CLK _14418_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15398_ hold517/A _15398_/CLK _15398_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13744__861 VPWR VGND VPWR VGND _15116_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_14349_ _14349_/Q _14349_/CLK _14349_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold605 hold605/X hold605/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 hold616/X hold616/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 hold627/X hold627/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 hold649/X hold649/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/X hold638/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09890_ VPWR VGND VGND VPWR _09890_/A _15480_/Q _09891_/S sky130_fd_sc_hd__nor2_1
XFILLER_69_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08910_ VPWR VGND VGND VPWR _08910_/X _15137_/Q _08924_/B sky130_fd_sc_hd__or2_1
X_08841_ VGND VPWR VPWR VGND _15172_/D fanout7/A _08842_/S hold812/X sky130_fd_sc_hd__mux2_1
Xhold1305 hold1305/X _14807_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 _10023_/A _15625_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1327 hold1327/X _15351_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1338 _09523_/A _14538_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08772_ VGND VPWR VPWR VGND _15234_/D _09860_/A0 _08772_/S hold265/X sky130_fd_sc_hd__mux2_1
Xhold1349 _09801_/A _14250_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07723_ VPWR VGND VPWR VGND _07827_/D _15587_/Q _07714_/X _07725_/B sky130_fd_sc_hd__a21o_1
X_07654_ VPWR VGND VGND VPWR _07857_/A _07654_/Y _07654_/B sky130_fd_sc_hd__nand2_1
X_07585_ VPWR VGND VGND VPWR _09010_/B _07586_/C _07585_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09324_ VGND VPWR VPWR VGND _09342_/S hold1092/X fanout49/X _14720_/D sky130_fd_sc_hd__mux2_2
X_13928__1045 VPWR VGND VPWR VGND _15300_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_09255_ VGND VPWR VPWR VGND _14788_/D fanout46/X _09269_/S hold706/X sky130_fd_sc_hd__mux2_1
X_08206_ VGND VPWR VGND VPWR _08206_/X _08280_/A2 _08203_/X _08201_/A _08205_/X sky130_fd_sc_hd__a211o_1
X_12959__76 VPWR VGND VPWR VGND _14202_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
Xclone49 VPWR VGND clone49/X clone49/A VPWR VGND sky130_fd_sc_hd__buf_6
X_09186_ VGND VPWR VPWR VGND _14905_/D hold322/X _09197_/S fanout12/X sky130_fd_sc_hd__mux2_1
X_08137_ VGND VPWR _08138_/B _08137_/B _08137_/A _08137_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_08068_ VPWR VGND VPWR VGND _15077_/Q _11440_/B _08068_/X _08293_/A3 _08041_/A _08067_/Y
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_1363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10030_ VGND VPWR VPWR VGND _10030_/A _15628_/D _10031_/C sky130_fd_sc_hd__xor2_1
X_11981_ VGND VPWR VPWR VGND _11981_/X _11978_/X _11995_/S _11977_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10932_ VPWR VGND VPWR VGND _10931_/X _11247_/A _12750_/B1 _10932_/X sky130_fd_sc_hd__a21o_1
X_10863_ VPWR VGND VGND VPWR _10863_/X hold630/A _10885_/S sky130_fd_sc_hd__or2_1
X_13687__804 VPWR VGND VPWR VGND _15027_/CLK clkload38/A sky130_fd_sc_hd__inv_2
XFILLER_73_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12602_ VPWR VGND VPWR VGND _12601_/X _12584_/A _12602_/B1 _12602_/X sky130_fd_sc_hd__a21o_1
X_10794_ VGND VPWR VPWR VGND _10794_/X _14206_/Q _10795_/S hold172/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15321_ _15321_/Q _15321_/CLK _15321_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12533_ VGND VPWR VPWR VGND _12533_/X hold695/A _12539_/S hold389/A sky130_fd_sc_hd__mux2_1
XFILLER_33_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13728__845 VPWR VGND VPWR VGND _15100_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_15252_ hold289/A _15252_/CLK _15252_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14203_ _14203_/Q _14203_/CLK _14203_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12464_ VGND VPWR VPWR VGND _12468_/B hold661/A _12479_/S hold223/A sky130_fd_sc_hd__mux2_1
X_11415_ VPWR VGND VGND VPWR _11415_/X _14821_/Q _14859_/Q sky130_fd_sc_hd__or2_1
X_15183_ hold501/A _15183_/CLK _15183_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1075 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12395_ VGND VPWR VGND VPWR _12395_/X _12720_/A1 _12391_/X _12394_/X _12485_/C1 sky130_fd_sc_hd__o211a_1
X_11346_ VPWR VGND VPWR VGND _11421_/A _11303_/A _14834_/Q _11347_/C _11313_/C sky130_fd_sc_hd__a22o_1
X_14134_ _14134_/Q _14134_/CLK _14134_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_4_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_10_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12973__90 VPWR VGND VPWR VGND _14216_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_11277_ VPWR VGND VGND VPWR _11561_/B _15440_/Q _11277_/B sky130_fd_sc_hd__or2_1
XFILLER_45_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10228_ VPWR VGND _10228_/X _10227_/X _10223_/X _10987_/S _10219_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10159_ VGND VPWR VPWR VGND _10159_/X _10158_/X _10467_/S _10157_/X sky130_fd_sc_hd__mux2_1
X_13280__397 VPWR VGND VPWR VGND _14555_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_14967_ hold532/A _14967_/CLK _14967_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14898_ hold578/A _14898_/CLK _14898_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_23_707 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_50_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07370_ VPWR VGND VGND VPWR _08201_/A _08201_/B _07369_/X _08180_/B sky130_fd_sc_hd__o21a_1
X_15519_ hold235/A _15519_/CLK _15519_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_751 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13174__291 VPWR VGND VPWR VGND _14449_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_09040_ VGND VPWR VPWR VGND _15050_/D hold663/X _09053_/S fanout41/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold402 hold402/X hold402/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 hold435/X hold435/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold413/X hold413/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 hold424/X hold424/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ VPWR VGND VGND VPWR _09942_/A _09943_/B _14130_/Q sky130_fd_sc_hd__nand2_1
Xhold468 hold468/X hold468/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 hold457/X hold457/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 hold446/X hold446/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold479 hold479/X hold479/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09873_ VPWR VGND VGND VPWR _09873_/A _09888_/S _09882_/A sky130_fd_sc_hd__nor2_1
X_13521__638 VPWR VGND VPWR VGND _14796_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
Xhold1124 hold1124/X _14240_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 hold1113/X _15417_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ VGND VPWR VPWR VGND _15189_/D fanout68/X _08846_/S hold737/X sky130_fd_sc_hd__mux2_1
XFILLER_6_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1102 hold1102/X _14877_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1157 hold1157/X _14302_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 hold1146/X _15223_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ VGND VPWR VPWR VGND _15251_/D fanout61/X _08776_/S hold313/X sky130_fd_sc_hd__mux2_1
Xhold1135 hold1135/X _15010_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1168 hold1168/X _14752_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 hold1179/X _15147_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07706_ VPWR VGND VGND VPWR _15565_/Q _07867_/B _07706_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08686_ VGND VPWR VGND VPWR _15286_/D hold950/X _08686_/A2 _08685_/X _12085_/C1 sky130_fd_sc_hd__o211a_1
X_07637_ VPWR VGND VGND VPWR _07637_/A _07637_/B _07637_/Y sky130_fd_sc_hd__nor2_1
X_07568_ VGND VPWR VPWR VGND _07568_/X _07558_/A _08880_/A _07567_/B _07567_/Y sky130_fd_sc_hd__o31a_4
X_13415__532 VPWR VGND VPWR VGND _14690_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_09307_ VGND VPWR VPWR VGND _14734_/D _09622_/A1 _09307_/S hold423/X sky130_fd_sc_hd__mux2_1
X_07499_ VGND VPWR VGND VPWR _07444_/X _08566_/B _07498_/X _07551_/B sky130_fd_sc_hd__o21bai_4
X_09238_ VPWR VGND VPWR VGND _08416_/Y _08415_/Y _09239_/B _14806_/D sky130_fd_sc_hd__a21oi_1
X_09169_ VGND VPWR VPWR VGND _14922_/D hold540/X _09191_/S clone146/X sky130_fd_sc_hd__mux2_1
X_12180_ VGND VPWR VPWR VGND _12180_/X _12179_/X _12180_/S _12178_/X sky130_fd_sc_hd__mux2_1
X_11200_ VPWR VGND VPWR VGND _11199_/X _11218_/A1 _11198_/X _11200_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11131_ VPWR VGND VGND VPWR _11131_/X _11143_/S _11131_/B sky130_fd_sc_hd__or2_1
Xhold980 hold980/X hold980/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 hold991/X hold991/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ VPWR VGND VGND VPWR _11247_/A _11062_/B _11062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_1205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10013_ VPWR VGND _10017_/C _10014_/B _15621_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_27_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14821_ _14821_/Q _14821_/CLK _14821_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_28_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14752_ _14752_/Q _14752_/CLK _14752_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11964_ VGND VPWR VPWR VGND _11964_/X _15491_/Q _11964_/S hold180/A sky130_fd_sc_hd__mux2_1
X_11895_ VPWR VGND VPWR VGND _11894_/X _11892_/X _11893_/X _11895_/X _12185_/A1 sky130_fd_sc_hd__a22o_1
XFILLER_45_887 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14683_ hold536/A _14683_/CLK _14683_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10915_ VPWR VGND VGND VPWR _10915_/X hold590/A _10924_/B sky130_fd_sc_hd__or2_1
X_10846_ VPWR VGND VPWR VGND _10843_/X _10846_/A1 _10845_/X _10846_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_879 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13158__275 VPWR VGND VPWR VGND _14433_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_15304_ _15304_/Q _15304_/CLK _15304_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10777_ VGND VPWR VGND VPWR _10777_/X hold979/A _11262_/A2 _10776_/X _10315_/S sky130_fd_sc_hd__o211a_1
XFILLER_13_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12516_ VGND VPWR VPWR VGND _12516_/X _14887_/Q _12664_/S hold371/A sky130_fd_sc_hd__mux2_1
X_15235_ hold161/A _15235_/CLK _15235_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12447_ VGND VPWR VGND VPWR _12447_/X _15022_/Q _12743_/A2 _12624_/S _12446_/X sky130_fd_sc_hd__o211a_1
X_15166_ hold842/A _15166_/CLK _15166_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12378_ VPWR VGND _12378_/X _12352_/X _12348_/X _12864_/A1 _12473_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_11329_ VGND VPWR VGND VPWR _14828_/D _07108_/Y _11327_/C _11328_/X _11327_/A sky130_fd_sc_hd__o211a_1
X_15097_ hold928/A _15097_/CLK _15097_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13927__1044 VPWR VGND VPWR VGND _15299_/CLK clkload15/A sky130_fd_sc_hd__inv_2
X_13856__973 VPWR VGND VPWR VGND _15228_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_36_821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08540_ VPWR VGND VPWR VGND _08540_/B1 _15315_/Q _08540_/A2 _08541_/B hold1420/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_640 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08471_ VGND VPWR VGND VPWR _08471_/X hold1242/X _08483_/A2 _08470_/X _09024_/A sky130_fd_sc_hd__o211a_1
XFILLER_63_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_36_865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07422_ VGND VPWR _07422_/X _08286_/A _15584_/Q _08286_/B VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_1_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07353_ _08006_/B _07267_/B _15459_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_17_1335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07284_ _07811_/A _07971_/A _07981_/A _07981_/B _07283_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_12929__46 VPWR VGND VPWR VGND _14172_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_17_Left_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09023_ VPWR VGND VPWR VGND _09022_/Y _09024_/A _09974_/A _15064_/D sky130_fd_sc_hd__a21oi_1
Xhold210 hold210/X hold210/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/X hold243/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/X hold221/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/X hold232/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold254/X hold254/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/X hold265/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/X hold287/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 hold276/X hold276/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ VPWR VGND VGND VPWR _09931_/C _09925_/Y _09925_/B sky130_fd_sc_hd__nand2_1
Xfanout701 VGND VPWR _12877_/S _12870_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout723 VGND VPWR _12750_/B1 _12713_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout712 VGND VPWR _08684_/S _08690_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold298 hold298/X hold298/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout734 VPWR VGND _12380_/B _11117_/B VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout756 VPWR VGND _07993_/A _07703_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout767 VGND VPWR _07420_/X _08293_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout745 VPWR VGND _08664_/B _08232_/B VPWR VGND sky130_fd_sc_hd__buf_2
X_09856_ VGND VPWR VPWR VGND _14166_/D hold651/X _09867_/S fanout14/X sky130_fd_sc_hd__mux2_1
Xfanout789 VPWR VGND _09890_/A _15478_/Q VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout778 VPWR VGND _08225_/C1 _07332_/Y VPWR VGND sky130_fd_sc_hd__buf_2
X_08807_ VGND VPWR VPWR VGND _15202_/D _09826_/A1 _08814_/S hold225/X sky130_fd_sc_hd__mux2_1
XFILLER_45_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09787_ VGND VPWR VPWR VGND _14262_/D fanout12/X _09798_/S hold459/X sky130_fd_sc_hd__mux2_1
XANTENNA_116 _09864_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08738_ VPWR VGND _14764_/D _08738_/B _14766_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XANTENNA_105 fanout424/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_54_651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_53_150 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08669_ VGND VPWR VPWR VGND _08669_/X _14402_/Q _08684_/S _14386_/Q sky130_fd_sc_hd__mux2_1
XFILLER_27_887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_27_876 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10700_ VGND VPWR VPWR VGND _10700_/X _15015_/Q _10700_/S hold419/A sky130_fd_sc_hd__mux2_1
XFILLER_14_526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_537 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11680_ VGND VPWR VPWR VGND _11680_/X hold863/A _12052_/S hold439/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10631_ VGND VPWR VPWR VGND _10631_/X hold407/A _10632_/B hold736/A sky130_fd_sc_hd__mux2_1
X_10562_ VPWR VGND VGND VPWR _10562_/X _14391_/Q _10562_/B sky130_fd_sc_hd__or2_1
X_12301_ VPWR VGND VGND VPWR _12301_/X hold209/A _12708_/S sky130_fd_sc_hd__or2_1
X_15020_ _15020_/Q _15020_/CLK _15020_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13799__916 VPWR VGND VPWR VGND _15171_/CLK clkload19/A sky130_fd_sc_hd__inv_2
X_10493_ VGND VPWR VPWR VGND _10493_/X hold822/A _10521_/B hold668/A sky130_fd_sc_hd__mux2_1
X_12232_ VPWR VGND VPWR VGND _12231_/X _12214_/A _11973_/B _12232_/X sky130_fd_sc_hd__a21o_1
X_12943__60 VPWR VGND VPWR VGND _14186_/CLK clkload44/A sky130_fd_sc_hd__inv_2
X_12163_ VGND VPWR VPWR VGND _12163_/X hold613/A _12171_/S hold442/A sky130_fd_sc_hd__mux2_1
X_13543__660 VPWR VGND VPWR VGND _14874_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_11114_ VPWR VGND VGND VPWR _11111_/X _11113_/X _10765_/S _11114_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12094_ VGND VPWR VPWR VGND _12098_/B hold384/A _12094_/S hold184/A sky130_fd_sc_hd__mux2_1
XFILLER_42_1417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11045_ VGND VPWR VPWR VGND _11049_/B hold889/A _11165_/S hold365/A sky130_fd_sc_hd__mux2_1
X_14122__1239 VPWR VGND VPWR VGND _15541_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_14804_ _14804_/Q clkload31/A _14804_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11947_ VGND VPWR VPWR VGND _11947_/X hold596/A _11950_/B hold304/A sky130_fd_sc_hd__mux2_1
XFILLER_29_191 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14735_ hold281/A _14735_/CLK _14735_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_632 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_835 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11878_ VGND VPWR VGND VPWR _11878_/X _11875_/X _11877_/X _11958_/A _12175_/A1 sky130_fd_sc_hd__a211o_1
X_14666_ _14666_/Q _14666_/CLK _14666_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10829_ VGND VPWR VGND VPWR _10829_/X _10828_/X _10827_/X _11205_/A _11104_/B1 sky130_fd_sc_hd__a211o_1
X_14597_ hold389/A _14597_/CLK _14597_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_20_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15218_ hold174/A _15218_/CLK _15218_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15149_ _15149_/Q _15149_/CLK _15149_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07971_ VPWR VGND VGND VPWR _07971_/A _10075_/A _07971_/Y sky130_fd_sc_hd__nor2_1
X_09710_ VGND VPWR VPWR VGND _14333_/D fanout39/X _09710_/S hold690/X sky130_fd_sc_hd__mux2_1
XFILLER_68_765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09641_ VGND VPWR VPWR VGND _14429_/D hold947/X _09656_/S fanout39/X sky130_fd_sc_hd__mux2_1
X_13592__709 VPWR VGND VPWR VGND _14923_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_09572_ VGND VPWR VPWR VGND _14493_/D hold1010/X _09584_/S fanout39/X sky130_fd_sc_hd__mux2_1
X_08523_ _08523_/X _15323_/Q _08523_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_71_919 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08454_ VPWR VGND VGND VPWR _08454_/X _15349_/Q _08488_/B sky130_fd_sc_hd__or2_1
XFILLER_51_687 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07405_ VPWR VGND _07637_/A _07636_/B _07639_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08385_ VGND VPWR VPWR VGND _15392_/D fanout71/X _08405_/S hold698/X sky130_fd_sc_hd__mux2_1
X_13486__603 VPWR VGND VPWR VGND _14761_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_07336_ _07621_/B _07162_/B _15473_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_09006_ VGND VPWR VGND VPWR _15102_/D hold1076/X _09015_/A2 _09005_/X _11337_/C1
+ sky130_fd_sc_hd__o211a_1
X_07267_ VPWR VGND VGND VPWR _15459_/Q _07267_/B _08028_/A sky130_fd_sc_hd__nor2_1
X_13527__644 VPWR VGND VPWR VGND _14807_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_07198_ VGND VPWR VPWR VGND _07376_/B _15599_/Q _07230_/S _14388_/Q sky130_fd_sc_hd__mux2_1
Xfanout531 VGND VPWR fanout538/X _12594_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout542 VGND VPWR _08491_/X _08522_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout520 VPWR VGND _12671_/S _12446_/B VPWR VGND sky130_fd_sc_hd__buf_2
X_09908_ _09909_/B _14766_/Q _09912_/A _14763_/Q _08507_/C _08529_/A VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__o311a_1
Xfanout564 _09637_/S _09656_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout553 VGND VPWR _08491_/A _07557_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout575 VPWR VGND _09377_/S _09346_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout586 VPWR VGND _09059_/S _09051_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09839_ VGND VPWR VPWR VGND _14183_/D hold643/X _09861_/S fanout78/X sky130_fd_sc_hd__mux2_1
Xfanout597 VPWR VGND _08806_/S _08780_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_12850_ VGND VPWR VPWR VGND _15574_/D _08216_/X _12860_/S _15574_/Q sky130_fd_sc_hd__mux2_1
XFILLER_41_1450 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11801_ VGND VPWR VPWR VGND _11801_/X hold862/A _12589_/S hold163/A sky130_fd_sc_hd__mux2_1
X_12781_ VPWR VGND VGND VPWR _12781_/A _12788_/S _12781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14520_ hold155/A _14520_/CLK _14520_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_42_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11732_ VGND VPWR VPWR VGND _11733_/B _11731_/Y _12472_/S _11723_/Y sky130_fd_sc_hd__mux2_1
X_11663_ VPWR VGND VGND VPWR _11663_/X hold649/A _11964_/S sky130_fd_sc_hd__or2_1
X_14451_ hold569/A _14451_/CLK _14451_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13926__1043 VPWR VGND VPWR VGND _15298_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_10614_ VGND VPWR VGND VPWR _10614_/X _10614_/A1 _10610_/X _10613_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
X_14382_ VGND VPWR VGND VPWR _14382_/Q _14382_/D clkload37/A sky130_fd_sc_hd__dfxtp_4
X_14200__918 _14200_/D _14200__918/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_11594_ VGND VPWR VPWR VGND _11594_/X hold626/A _11756_/S hold892/A sky130_fd_sc_hd__mux2_1
X_10545_ VPWR VGND VPWR VGND _10544_/X _10662_/S _10667_/C1 _10545_/X sky130_fd_sc_hd__a21o_1
X_10476_ VGND VPWR VPWR VGND _10476_/X hold781/A _10484_/B hold699/A sky130_fd_sc_hd__mux2_1
X_12215_ VPWR VGND VGND VPWR _12215_/X hold591/A _12220_/S sky130_fd_sc_hd__or2_1
X_15003_ _15003_/Q _15003_/CLK _15003_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12146_ VGND VPWR VPWR VGND _12146_/X hold918/A _12205_/S hold723/A sky130_fd_sc_hd__mux2_1
XFILLER_69_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12077_ VGND VPWR VGND VPWR _12077_/X _15012_/Q _12229_/A2 _12069_/S _12076_/X sky130_fd_sc_hd__o211a_1
X_11028_ VGND VPWR VPWR VGND _11028_/X hold845/A _11175_/S hold386/A sky130_fd_sc_hd__mux2_1
X_13320__437 VPWR VGND VPWR VGND _14595_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_15698_ VPWR VGND uo_out[3] _15698_/A VPWR VGND sky130_fd_sc_hd__buf_2
X_14718_ hold762/A _14718_/CLK _14718_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Left_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14649_ hold667/A _14649_/CLK _14649_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08170_ VGND VPWR VGND VPWR _08170_/X _08299_/A2 _08152_/X _15613_/Q _08169_/X sky130_fd_sc_hd__a211o_1
XANTENNA_27 _14404_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_16 _09557_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_38 _12864_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07121_ VPWR VGND VPWR VGND _09970_/A _15162_/Q sky130_fd_sc_hd__inv_2
XANTENNA_49 _08178_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_13214__331 VPWR VGND VPWR VGND _14489_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XFILLER_9_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_34_Left_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07954_ VGND VPWR VPWR VGND _15531_/D _07953_/X _07954_/S hold206/X sky130_fd_sc_hd__mux2_1
XFILLER_25_1445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07885_ VPWR VGND VGND VPWR _07885_/A _07886_/B _07885_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09624_ VGND VPWR VPWR VGND _14444_/D fanout98/X _09625_/S hold520/X sky130_fd_sc_hd__mux2_1
XFILLER_44_919 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09555_ VGND VPWR VPWR VGND _14507_/D _08299_/X _09555_/S hold214/X sky130_fd_sc_hd__mux2_1
X_08506_ VPWR VGND VPWR VGND _09909_/A _08508_/B sky130_fd_sc_hd__inv_2
X_09486_ _09486_/B _09486_/X _09486_/A _09486_/C VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_43_Left_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08437_ VGND VPWR VGND VPWR _15358_/D _15357_/Q _08448_/B _08436_/X _11382_/S sky130_fd_sc_hd__o211a_1
X_14121__1238 VPWR VGND VPWR VGND _15540_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_08368_ VGND VPWR VPWR VGND _15405_/D hold818/X _08375_/S _09860_/A0 sky130_fd_sc_hd__mux2_1
X_08299_ VGND VPWR VGND VPWR _08299_/X _08299_/A2 hold807/A _08294_/X _08298_/X sky130_fd_sc_hd__a211o_2
X_07319_ VPWR VGND VGND VPWR _15471_/Q _07319_/B _07339_/B sky130_fd_sc_hd__nor2_1
X_10330_ VGND VPWR VPWR VGND _10330_/X _15005_/Q _11102_/S hold759/A sky130_fd_sc_hd__mux2_1
X_13761__878 VPWR VGND VPWR VGND _15133_/CLK clkload19/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_52_Left_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10261_ VGND VPWR VPWR VGND _10261_/X hold609/A _11240_/S hold768/A sky130_fd_sc_hd__mux2_1
XFILLER_79_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12000_ VGND VPWR VGND VPWR _12000_/X _12008_/C1 _11995_/X _11999_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
X_10192_ VPWR VGND VGND VPWR _10192_/X _14381_/Q _10192_/B sky130_fd_sc_hd__or2_1
X_12913__30 VPWR VGND VPWR VGND _14156_/CLK clkload7/A sky130_fd_sc_hd__inv_2
Xfanout350 VGND VPWR _10144_/S _10613_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout372 VPWR VGND _11250_/S fanout381/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout361 VPWR VGND _10662_/S _08195_/C VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout383 VGND VPWR fanout390/X _10614_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1005 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_59_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout394 VGND VPWR _10890_/A _11004_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_74_565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_1280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13655__772 VPWR VGND VPWR VGND _14995_/CLK clkload38/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_61_Left_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12833_ VGND VPWR VPWR VGND _12833_/B _07846_/B _12833_/A _12833_/X sky130_fd_sc_hd__or3b_1
X_15621_ _15621_/Q clkload50/A _15621_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15552_ _15552_/Q clkload31/A _15552_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12764_ VGND VPWR VPWR VGND _12765_/B _08186_/Y _12820_/B _08187_/Y sky130_fd_sc_hd__mux2_1
X_15483_ hold809/A _15483_/CLK _15483_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14503_ hold751/A _14503_/CLK _14503_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11715_ VPWR VGND VGND VPWR _11696_/Y _11714_/X _12380_/B _15448_/Q _15448_/D _12085_/C1
+ sky130_fd_sc_hd__o221a_1
X_12695_ VPWR VGND VGND VPWR _12732_/A _12695_/B _12695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11646_ VPWR VGND VGND VPWR _11646_/X _11948_/S _11646_/B sky130_fd_sc_hd__or2_1
X_14434_ hold774/A _14434_/CLK _14434_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14365_ hold869/A _14365_/CLK _14365_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11577_ VGND VPWR VPWR VGND _11577_/X hold366/A _12086_/S hold563/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Left_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold809 hold809/X hold809/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10528_ VGND VPWR VPWR VGND _10528_/X hold763/A _10627_/S hold848/A sky130_fd_sc_hd__mux2_1
X_14296_ hold514/A _14296_/CLK _14296_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10459_ VGND VPWR VPWR VGND _10459_/X _10456_/X _10467_/S _10455_/X sky130_fd_sc_hd__mux2_1
X_12129_ VGND VPWR VPWR VGND _12129_/X _12126_/X _12147_/S _12125_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07670_ VGND VPWR VGND VPWR _07670_/X _07665_/A _07859_/B _07668_/Y _07669_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09340_ VGND VPWR VPWR VGND _14704_/D hold494/X _09345_/S _09688_/A0 sky130_fd_sc_hd__mux2_1
X_09271_ VGND VPWR VPWR VGND _14772_/D _09829_/A1 _09272_/S hold753/X sky130_fd_sc_hd__mux2_1
X_08222_ VGND VPWR VPWR VGND _08223_/A _08222_/X _08222_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08153_ VGND VPWR VPWR VGND _08153_/A _08153_/X _08153_/B sky130_fd_sc_hd__xor2_1
X_07104_ VPWR VGND VPWR VGND _08902_/A _15141_/Q sky130_fd_sc_hd__inv_2
X_08084_ VPWR VGND VGND VPWR _08277_/S _10063_/A _08084_/Y sky130_fd_sc_hd__nor2_1
X_13598__715 VPWR VGND VPWR VGND _14938_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_08986_ VPWR VGND VGND VPWR _09007_/A _08986_/B _08986_/Y sky130_fd_sc_hd__nor2_1
X_07937_ VPWR VGND VPWR VGND _12472_/S _08286_/A clone17/A _07953_/A sky130_fd_sc_hd__a21oi_1
XFILLER_29_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_56_521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13639__756 VPWR VGND VPWR VGND _14979_/CLK clkload14/A sky130_fd_sc_hd__inv_2
X_13925__1042 VPWR VGND VPWR VGND _15297_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_07868_ VGND VPWR VPWR VGND _07868_/A _07869_/B _07868_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_779 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09607_ VGND VPWR VPWR VGND _14461_/D fanout40/X _09622_/S hold867/X sky130_fd_sc_hd__mux2_1
X_07799_ _07800_/B _07958_/B _07958_/C _07958_/D _07958_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_43_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09538_ VGND VPWR VPWR VGND _14524_/D fanout37/X _09553_/S hold316/X sky130_fd_sc_hd__mux2_1
X_09469_ VGND VPWR VPWR VGND _14587_/D fanout32/X _09485_/S hold442/X sky130_fd_sc_hd__mux2_1
X_11500_ VGND VPWR VPWR VGND _11500_/X _11499_/X _11537_/S _15464_/Q sky130_fd_sc_hd__mux2_1
X_12480_ VGND VPWR VGND VPWR _12480_/X _12479_/X _12478_/X _12476_/S _12485_/C1 sky130_fd_sc_hd__a211o_1
X_11431_ VGND VPWR VGND VPWR _14930_/D hold1408/X _11431_/A2 _11430_/X _11431_/C1
+ sky130_fd_sc_hd__o211a_1
X_14150_ _14150_/Q _14150_/CLK _14150_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11362_ _11362_/X _14859_/Q _14821_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_10313_ VGND VPWR VPWR VGND _10313_/X _14193_/Q _11098_/S hold243/A sky130_fd_sc_hd__mux2_1
X_11293_ VGND VPWR VPWR VGND _11294_/B _14815_/Q _11299_/S _14383_/Q sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_5_Left_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10244_ VGND VPWR VGND VPWR _10244_/X _11235_/A1 _10240_/X _10243_/X _10918_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_3_366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10175_ VPWR VGND VPWR VGND _10174_/X _10703_/A _10706_/C1 _10175_/X sky130_fd_sc_hd__a21o_1
Xfanout191 VGND VPWR _12684_/S _12698_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_14983_ hold419/A _14983_/CLK _14983_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout180 VPWR VGND _12470_/S _12367_/S VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_35_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13391__508 VPWR VGND VPWR VGND _14666_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_12816_ VGND VPWR VPWR VGND _12817_/B _07931_/X _12820_/B _07915_/Y sky130_fd_sc_hd__mux2_1
X_15604_ _15604_/Q clkload19/A _15604_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14206__924 _14206_/D _14206__924/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_13432__549 VPWR VGND VPWR VGND _14707_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_12747_ VGND VPWR VPWR VGND _12747_/X _15397_/Q _12747_/S _15544_/Q sky130_fd_sc_hd__mux2_1
X_15535_ hold288/A _15535_/CLK _15535_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15466_ _15466_/Q clkload45/A _15466_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12678_ VGND VPWR VPWR VGND _12682_/B hold500/A _12701_/S hold577/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14417_ hold962/A _14417_/CLK _14417_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11629_ VGND VPWR VGND VPWR _11629_/X _11628_/X _11627_/X _11625_/S _12099_/C1 sky130_fd_sc_hd__a211o_1
X_15397_ _15397_/Q _15397_/CLK _15397_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold606 hold606/X hold606/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13285__402 VPWR VGND VPWR VGND _14560_/CLK clkload48/A sky130_fd_sc_hd__inv_2
Xhold617 hold617/X hold617/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14348_ hold871/A _14348_/CLK _14348_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold639 hold639/X hold639/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 hold628/X hold628/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ _14279_/Q _14279_/CLK _14279_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08840_ VGND VPWR VPWR VGND _15173_/D fanout9/A _08850_/S hold794/X sky130_fd_sc_hd__mux2_1
XFILLER_58_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13326__443 VPWR VGND VPWR VGND _14601_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
XFILLER_58_819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1306 hold1306/X _14847_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 hold1339/X _15141_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1328 hold1328/X _15133_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08771_ VGND VPWR VPWR VGND _15235_/D _09859_/A0 _08779_/S hold161/X sky130_fd_sc_hd__mux2_1
Xhold1317 hold1317/X _15065_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14120__1237 VPWR VGND VPWR VGND _15539_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_07722_ VPWR VGND VPWR VGND _07722_/Y _07938_/B sky130_fd_sc_hd__inv_2
XFILLER_38_598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07653_ VGND VPWR _07654_/B _07653_/A _07653_/B VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07584_ VPWR VGND VPWR VGND _07585_/B _07587_/B sky130_fd_sc_hd__inv_2
XFILLER_55_1202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09323_ VGND VPWR VPWR VGND _14721_/D hold465/X _09327_/S clone5/A sky130_fd_sc_hd__mux2_1
X_09254_ VGND VPWR VPWR VGND _09272_/S fanout48/X hold1189/X _14789_/D sky130_fd_sc_hd__mux2_2
Xclone17 VPWR VGND clone17/X clone17/A VPWR VGND sky130_fd_sc_hd__buf_6
X_08205_ VPWR VGND VPWR VGND _15070_/Q _08293_/B1 _08205_/X _08263_/A2 _07213_/X _08204_/X
+ sky130_fd_sc_hd__a221o_1
X_09185_ VGND VPWR VPWR VGND _14906_/D hold858/X _09197_/S fanout15/X sky130_fd_sc_hd__mux2_1
X_08136_ VPWR VGND VGND VPWR _08136_/A _08136_/B _12774_/B sky130_fd_sc_hd__nor2_1
X_08067_ VPWR VGND VGND VPWR _08067_/A _08104_/B _08067_/Y sky130_fd_sc_hd__nor2_1
X_13069__186 VPWR VGND VPWR VGND _14312_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_08969_ VPWR VGND VGND VPWR _08969_/X _08969_/A _08969_/B sky130_fd_sc_hd__or2_1
X_11980_ VGND VPWR VGND VPWR _11980_/X _12008_/A1 _11976_/X _11979_/X _12017_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_5_1199 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10931_ VPWR VGND _10931_/X _10930_/X _10926_/X _10987_/S _10922_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10862_ VGND VPWR VPWR VGND _10862_/X _10861_/X _11110_/A _10860_/X sky130_fd_sc_hd__mux2_1
X_12601_ VPWR VGND _12601_/X _12600_/X _12596_/X _12583_/S _12592_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10793_ VGND VPWR VGND VPWR _10793_/X _11218_/A1 _10788_/X _10792_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_31_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15320_ _15320_/Q _15320_/CLK _15320_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12532_ VGND VPWR VPWR VGND _12532_/X hold946/A _12539_/S hold893/A sky130_fd_sc_hd__mux2_1
X_13767__884 VPWR VGND VPWR VGND _15139_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_15251_ hold313/A _15251_/CLK _15251_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12463_ VPWR VGND VPWR VGND _12462_/X _12722_/A1 _12461_/X _12463_/Y sky130_fd_sc_hd__a21oi_1
X_11414_ VGND VPWR VGND VPWR _14858_/D _07106_/Y _11411_/X _11413_/X _08541_/A sky130_fd_sc_hd__o211a_1
X_14202_ _14202_/Q _14202_/CLK _14202_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15182_ hold853/A _15182_/CLK _15182_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12394_ VPWR VGND VGND VPWR _12394_/X _12396_/S _12394_/B sky130_fd_sc_hd__or2_1
X_11345_ VPWR VGND _14833_/D _11410_/A _14833_/Q _11327_/A _11344_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14133_ hold539/A _14133_/CLK _14133_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13013__130 VPWR VGND VPWR VGND _14256_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_11276_ VPWR VGND VGND VPWR _11277_/B _15439_/Q _11557_/B sky130_fd_sc_hd__or2_1
XFILLER_10_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10227_ VGND VPWR VGND VPWR _10227_/X _10224_/X _10226_/X _11004_/A1 _11237_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_45_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10158_ VGND VPWR VPWR VGND _10158_/X _14477_/Q _10169_/B hold636/A sky130_fd_sc_hd__mux2_1
XFILLER_66_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_43_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14966_ _14966_/Q _14966_/CLK _14966_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10089_ VGND VPWR VPWR VGND _10089_/X _10086_/X _10613_/A _10085_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_833 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14897_ hold499/A _14897_/CLK _14897_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15518_ hold314/A _15518_/CLK _15518_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13924__1041 VPWR VGND VPWR VGND _15296_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_15449_ _15449_/Q clkload35/A _15449_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
Xhold414 hold414/X hold414/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 hold436/X hold436/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 hold425/X hold425/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 hold403/X hold403/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ VPWR VGND VGND VPWR _09947_/C _14131_/Q _14130_/Q sky130_fd_sc_hd__or2_1
Xhold458 hold458/X hold458/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 hold447/X hold447/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 hold469/X hold469/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13560__677 VPWR VGND VPWR VGND _14891_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_09872_ VGND VPWR _09880_/B _09871_/Y _14152_/D _09906_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_08823_ VGND VPWR VPWR VGND _15190_/D fanout73/X _08846_/S hold691/X sky130_fd_sc_hd__mux2_1
Xhold1103 hold1103/X _15029_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 hold1114/X _15025_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 hold1125/X _15104_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1158 hold1158/X _14753_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1147 hold1147/X _14916_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 hold1136/X _14863_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ VGND VPWR VPWR VGND _15252_/D fanout65/X _08773_/S hold289/X sky130_fd_sc_hd__mux2_1
Xhold1169 _09940_/S _14131_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ VPWR VGND VGND VPWR _07867_/A _15565_/Q _07706_/B sky130_fd_sc_hd__or2_1
XFILLER_2_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08685_ VPWR VGND VPWR VGND _15285_/Q _08562_/A _08685_/X _08691_/B1 _08684_/X _08688_/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07636_ VPWR VGND VGND VPWR _07639_/A _07636_/B _07637_/B sky130_fd_sc_hd__nor2_1
X_07567_ VPWR VGND VGND VPWR _15347_/Q _07567_/Y _07567_/B sky130_fd_sc_hd__nand2_1
X_13454__571 VPWR VGND VPWR VGND _14729_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_41_549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_55_1043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09306_ VGND VPWR VPWR VGND _14735_/D _09829_/A1 _09307_/S hold281/X sky130_fd_sc_hd__mux2_1
X_09237_ VPWR VGND VGND VPWR _09237_/C _09237_/B _09239_/B _14807_/D sky130_fd_sc_hd__nor3_1
X_07498_ VPWR VGND VGND VPWR _07498_/X _07714_/A _15457_/Q _15458_/Q _15459_/Q _15460_/Q
+ sky130_fd_sc_hd__o41a_1
XFILLER_33_1363 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_1385 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_428 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09168_ VGND VPWR VPWR VGND _14923_/D hold424/X _09191_/S fanout80/X sky130_fd_sc_hd__mux2_1
X_08119_ VPWR VGND VGND VPWR _08119_/X _08277_/S _10063_/C sky130_fd_sc_hd__or2_1
X_09099_ VGND VPWR VPWR VGND _14996_/D hold340/X _09124_/S fanout80/X sky130_fd_sc_hd__mux2_1
X_13801__918 VPWR VGND VPWR VGND _15173_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_11130_ VGND VPWR VPWR VGND _11130_/X hold582/A _11142_/S hold287/A sky130_fd_sc_hd__mux2_1
Xhold970 hold970/X hold970/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/X hold981/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 hold992/X hold992/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ VGND VPWR VPWR VGND _11062_/B _11060_/Y _11246_/S _11052_/Y sky130_fd_sc_hd__mux2_1
XFILLER_49_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10012_ VPWR VGND VGND VPWR _10014_/B _10012_/B _15620_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14820_ _14820_/Q _14821_/CLK _14820_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14751_ hold217/A _14751_/CLK _14751_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11963_ VGND VPWR VPWR VGND _11963_/X _15009_/Q _11964_/S hold391/A sky130_fd_sc_hd__mux2_1
X_11894_ VGND VPWR VPWR VGND _11894_/X _11891_/X _11894_/S _11890_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14682_ hold558/A _14682_/CLK _14682_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10914_ VPWR VGND VGND VPWR _11247_/A _10914_/B _10914_/Y sky130_fd_sc_hd__nor2_1
X_10845_ VPWR VGND VPWR VGND _10844_/X _10315_/S _11259_/C1 _10845_/X sky130_fd_sc_hd__a21o_1
XFILLER_44_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15303_ hold986/A _15303_/CLK _15303_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10776_ VPWR VGND VGND VPWR _10776_/X hold685/A _10850_/S sky130_fd_sc_hd__or2_1
XFILLER_13_785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_51_1430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12515_ VGND VPWR VGND VPWR _12515_/X hold845/A _12669_/A2 _12662_/A1 _12514_/X sky130_fd_sc_hd__o211a_1
XFILLER_9_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15234_ hold265/A _15234_/CLK _15234_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12446_ VPWR VGND VGND VPWR _12446_/X hold471/A _12446_/B sky130_fd_sc_hd__or2_1
X_12377_ VGND VPWR VPWR VGND _12377_/X _12376_/X _12472_/S _12368_/X sky130_fd_sc_hd__mux2_1
X_15165_ hold984/A _15165_/CLK _15165_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11328_ VGND VPWR _14825_/Q _11313_/C _14826_/Q _11328_/X _14828_/Q _14827_/Q VPWR
+ VGND sky130_fd_sc_hd__a41o_1
X_15096_ _15096_/Q clkload37/A _15096_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_4_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_45_1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11259_ VGND VPWR VGND VPWR _11259_/X _11256_/X _11258_/X _10816_/A _11259_/C1 sky130_fd_sc_hd__a211o_1
X_13397__514 VPWR VGND VPWR VGND _14672_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
XFILLER_10_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_844 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14949_ hold801/A _14949_/CLK _14949_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08470_ VPWR VGND VGND VPWR _08470_/X _15341_/Q _08484_/B sky130_fd_sc_hd__or2_1
XFILLER_51_803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13438__555 VPWR VGND VPWR VGND _14713_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_07421_ VPWR VGND VGND VPWR _07421_/Y _07421_/A _08286_/B sky130_fd_sc_hd__nand2_2
X_07352_ VGND VPWR VGND VPWR _07263_/B _07982_/B _15460_/Q sky130_fd_sc_hd__nand2b_2
X_07283_ VPWR VGND VPWR VGND _07283_/Y _07916_/B _07286_/B _07279_/Y _07288_/A sky130_fd_sc_hd__a211oi_1
X_09022_ VPWR VGND VGND VPWR _15697_/A _09022_/B _09022_/Y sky130_fd_sc_hd__nor2_1
Xhold200 hold200/X hold200/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 hold211/X hold211/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/X hold244/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/X hold222/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/X hold233/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 hold277/X hold277/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/X hold255/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/X hold266/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ VPWR VGND _14140_/Q _14136_/Q _09923_/D _09925_/B _14135_/Q VPWR VGND sky130_fd_sc_hd__o31ai_1
Xfanout702 VPWR VGND _12877_/S _10054_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout713 VPWR VGND _08684_/S _08687_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout724 VPWR VGND _12750_/B1 _11974_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xhold288 hold288/X hold288/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 hold299/X hold299/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout757 VPWR VGND _10060_/C _08604_/B2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout735 VGND VPWR _09975_/Y _12807_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09855_ VGND VPWR VPWR VGND _14167_/D hold848/X _09867_/S fanout16/X sky130_fd_sc_hd__mux2_1
XFILLER_28_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout746 VGND VPWR _08640_/B _08232_/B VPWR VGND sky130_fd_sc_hd__buf_1
X_08806_ VGND VPWR VPWR VGND _15203_/D _09825_/A1 _08806_/S hold252/X sky130_fd_sc_hd__mux2_1
Xfanout768 VPWR VGND _10072_/B _07420_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout779 VPWR VGND _07304_/B1 _07265_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_39_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09786_ VGND VPWR VPWR VGND _14263_/D fanout17/X _09798_/S hold771/X sky130_fd_sc_hd__mux2_1
X_08737_ _08737_/X _15698_/A _09938_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XANTENNA_106 fanout424/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk _12923__40/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XANTENNA_117 _09126_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_38_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08668_ VGND VPWR VGND VPWR _15292_/D hold1025/X _08721_/A2 _08667_/X _11937_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_685 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07619_ VPWR VGND VGND VPWR _07163_/A _07619_/B _07620_/B sky130_fd_sc_hd__nand2b_1
XFILLER_74_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08599_ VGND VPWR VPWR VGND _08998_/B _15550_/Q _07552_/B1 _08604_/B2 _08598_/Y sky130_fd_sc_hd__o2bb2a_1
X_10630_ VGND VPWR VGND VPWR _10630_/X _10627_/X _10629_/X _10634_/A1 _10630_/C1 sky130_fd_sc_hd__a211o_1
X_13190__307 VPWR VGND VPWR VGND _14465_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_10561_ VPWR VGND VPWR VGND _10561_/X _10618_/A _10534_/X _10542_/X _10560_/X _10559_/X
+ sky130_fd_sc_hd__o32a_1
X_12300_ VGND VPWR VGND VPWR _12300_/X _12297_/X _12299_/X _12748_/A1 _12744_/C1 sky130_fd_sc_hd__a211o_1
X_13231__348 VPWR VGND VPWR VGND _14506_/CLK clkload44/A sky130_fd_sc_hd__inv_2
X_10492_ VGND VPWR VPWR VGND _10492_/X hold739/A _10521_/B hold232/A sky130_fd_sc_hd__mux2_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12231_ VPWR VGND _12231_/X _12230_/X _12226_/X _12139_/S _12222_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12162_ VGND VPWR VPWR VGND _12162_/X hold938/A _12171_/S hold231/A sky130_fd_sc_hd__mux2_1
X_11113_ VGND VPWR VGND VPWR _11113_/X _11110_/A _11109_/X _11112_/X _11263_/C1 sky130_fd_sc_hd__o211a_1
X_13084__201 VPWR VGND VPWR VGND _14327_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_13879__996 VPWR VGND VPWR VGND _15251_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_12093_ VPWR VGND VPWR VGND _12092_/X _12101_/A1 _12091_/X _12093_/Y sky130_fd_sc_hd__a21oi_1
X_11044_ VPWR VGND VGND VPWR _11025_/Y _11043_/X _12677_/A2 _14404_/Q _14404_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_13125__242 VPWR VGND VPWR VGND _14368_/CLK clkload48/A sky130_fd_sc_hd__inv_2
XFILLER_42_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14803_ _14803_/Q clkload31/A _14803_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13923__1040 VPWR VGND VPWR VGND _15295_/CLK clkload13/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_56_clk clkload35/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_75_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11946_ VGND VPWR VPWR VGND _11946_/X _14197_/Q _11950_/B hold478/A sky130_fd_sc_hd__mux2_1
X_14734_ hold423/A _14734_/CLK _14734_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11877_ VGND VPWR VGND VPWR _11877_/X hold951/A _12192_/A2 _12174_/S _11876_/X sky130_fd_sc_hd__o211a_1
X_14665_ hold577/A _14665_/CLK _14665_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10828_ VGND VPWR VPWR VGND _10828_/X hold571/A _11093_/S hold526/A sky130_fd_sc_hd__mux2_1
XFILLER_38_1071 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14596_ hold467/A _14596_/CLK _14596_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10759_ VGND VPWR VPWR VGND _10759_/X _14205_/Q _10835_/B hold277/A sky130_fd_sc_hd__mux2_1
X_15217_ _15217_/Q _15217_/CLK _15217_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13823__940 VPWR VGND VPWR VGND _15195_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XFILLER_58_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12989__106 VPWR VGND VPWR VGND _14232_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_12429_ VGND VPWR VPWR VGND _12429_/X _14210_/Q _12651_/S hold174/A sky130_fd_sc_hd__mux2_1
X_15148_ _15148_/Q _15148_/CLK _15148_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07970_ VGND VPWR VGND VPWR _07970_/X _07966_/A _10064_/A _07966_/Y _10071_/A sky130_fd_sc_hd__o211a_1
X_15079_ _15079_/Q clkload37/A _15079_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09640_ VGND VPWR VPWR VGND _14430_/D _09656_/S hold1235/X clone44/X sky130_fd_sc_hd__mux2_4
XFILLER_3_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09571_ VGND VPWR VPWR VGND _14494_/D _09587_/S hold1229/X fanout42/X sky130_fd_sc_hd__mux2_4
X_08522_ _08522_/X _08523_/B _08522_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_47_clk _12969__86/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_13672__789 VPWR VGND VPWR VGND _15012_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_08453_ VGND VPWR VGND VPWR _15350_/D _15349_/Q _08448_/B _08452_/X _11308_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_24_836 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07404_ VPWR VGND VGND VPWR _07665_/B _07403_/X _07343_/X _07636_/B sky130_fd_sc_hd__o21a_1
XFILLER_24_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08384_ VGND VPWR VPWR VGND _15393_/D _08393_/S fanout72/X hold1245/X sky130_fd_sc_hd__mux2_4
X_07335_ _07335_/X _07157_/B _15474_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_07266_ VPWR VGND _07268_/A _07267_/B _15459_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_09005_ VGND VPWR VGND VPWR _09005_/X _09007_/A _09016_/B1 hold971/X _09004_/Y sky130_fd_sc_hd__a211o_1
X_07197_ VPWR VGND VPWR VGND _07248_/A _07197_/A sky130_fd_sc_hd__inv_2
X_13566__683 VPWR VGND VPWR VGND _14897_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_09907_ VGND VPWR VPWR VGND _14141_/D hold819/X _09907_/S _09906_/Y sky130_fd_sc_hd__mux2_1
XFILLER_59_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout532 VGND VPWR _12282_/S _12701_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13109__226 VPWR VGND VPWR VGND _14352_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
Xfanout510 VGND VPWR _12409_/B _11748_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout521 VGND VPWR _12446_/B _12661_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout565 _09656_/S _09626_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout543 VPWR VGND VGND VPWR clone18/A _07873_/B1 sky130_fd_sc_hd__buf_12
Xfanout554 _09833_/S _09825_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_24_1115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout576 _09357_/S _09376_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout598 _08808_/S _08811_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_47_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09838_ VGND VPWR VPWR VGND _09861_/S hold1153/X clone49/X _14184_/D sky130_fd_sc_hd__mux2_2
Xfanout587 VGND VPWR _09026_/X _09051_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09769_ VGND VPWR VPWR VGND _14280_/D clone45/X _09792_/S hold535/X sky130_fd_sc_hd__mux2_1
X_11800_ VGND VPWR VPWR VGND _11800_/X _14193_/Q _12589_/S hold243/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_clk _12974__91/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12780_ VGND VPWR _08585_/Y _12779_/Y _15552_/D _10060_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_42_655 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11731_ VPWR VGND VPWR VGND _11730_/X _12415_/C1 _11729_/X _11731_/Y sky130_fd_sc_hd__a21oi_1
X_11662_ VGND VPWR VPWR VGND _11662_/X _11661_/X _12180_/S _11660_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14450_ _14450_/Q _14450_/CLK _14450_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_817 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14381_ VGND VPWR VGND VPWR _14381_/Q _14381_/D clkload23/A sky130_fd_sc_hd__dfxtp_4
X_11593_ VGND VPWR VGND VPWR _11593_/X _12101_/A1 _11588_/X _11592_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
X_10613_ VPWR VGND VGND VPWR _10613_/X _10613_/A _10613_/B sky130_fd_sc_hd__or2_1
X_13807__924 VPWR VGND VPWR VGND _15179_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_10544_ VGND VPWR VPWR VGND _10544_/X _14359_/Q _10554_/S hold502/A sky130_fd_sc_hd__mux2_1
X_10475_ VGND VPWR VGND VPWR _10475_/X hold830/A _10688_/A2 _10474_/X _10486_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_6_589 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12214_ VPWR VGND VGND VPWR _12214_/A _12214_/B _12214_/Y sky130_fd_sc_hd__nor2_1
X_15002_ _15002_/Q _15002_/CLK _15002_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12145_ VGND VPWR VPWR VGND _12145_/X hold874/A _12205_/S hold558/A sky130_fd_sc_hd__mux2_1
XFILLER_37_8 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12076_ VPWR VGND VGND VPWR _12076_/X hold335/A _12227_/S sky130_fd_sc_hd__or2_1
X_11027_ VGND VPWR VGND VPWR _11027_/X _14887_/Q _11184_/A2 _11026_/X _11176_/S sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_29_clk clkload46/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_15697_ VPWR VGND uo_out[2] _15697_/A VPWR VGND sky130_fd_sc_hd__buf_2
X_14717_ hold742/A _14717_/CLK _14717_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11929_ VGND VPWR VGND VPWR _11929_/X hold750/A _12229_/A2 _11925_/S _11928_/X sky130_fd_sc_hd__o211a_1
X_14648_ hold654/A _14648_/CLK _14648_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1420 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_39 _12213_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_28 _14404_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_17 _09591_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_07120_ VPWR VGND VPWR VGND _08500_/B _15365_/Q sky130_fd_sc_hd__inv_2
X_13253__370 VPWR VGND VPWR VGND _14528_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_14579_ hold178/A _14579_/CLK _14579_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13600__717 VPWR VGND VPWR VGND _14940_/CLK clkload11/A sky130_fd_sc_hd__inv_2
XFILLER_68_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07953_ VPWR VGND VPWR VGND _07953_/B _07953_/C _07953_/A _07953_/X sky130_fd_sc_hd__or3_4
X_07884_ VPWR VGND VGND VPWR _07885_/B _15564_/Q _07906_/A sky130_fd_sc_hd__or2_1
XFILLER_25_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09623_ VGND VPWR VPWR VGND _14445_/D _09865_/A0 _09625_/S hold681/X sky130_fd_sc_hd__mux2_1
XFILLER_58_1222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09554_ VGND VPWR VPWR VGND _14508_/D _09658_/A0 _09555_/S hold250/X sky130_fd_sc_hd__mux2_1
X_08505_ VPWR VGND VGND VPWR _08505_/C _09923_/D _08505_/A _08508_/B sky130_fd_sc_hd__nor3_1
X_09485_ VGND VPWR VPWR VGND _14571_/D fanout95/X _09485_/S hold199/X sky130_fd_sc_hd__mux2_1
X_08436_ VPWR VGND VGND VPWR _08436_/X _15358_/Q _08488_/B sky130_fd_sc_hd__or2_1
XFILLER_51_463 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08367_ VGND VPWR VPWR VGND _15406_/D hold725/X _08375_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
X_07318_ VGND VPWR VGND VPWR _07663_/B _07313_/B _07679_/A _07313_/A _07693_/B sky130_fd_sc_hd__a211o_1
XFILLER_32_1417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08298_ VGND VPWR VPWR VGND _08298_/X _10058_/A1 _08297_/X _08295_/Y _08172_/X _08298_/A1
+ sky130_fd_sc_hd__o2111a_1
X_07249_ VPWR VGND _08062_/A _07249_/B _07249_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_10260_ VGND VPWR VGND VPWR _10260_/X _10257_/X _10259_/X _11235_/A1 _10918_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_69_1384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10191_ VPWR VGND VPWR VGND _10191_/X _10507_/A _10164_/X _10172_/X _10190_/X _10189_/X
+ sky130_fd_sc_hd__o32a_1
Xfanout340 VGND VPWR _11107_/S _11098_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout351 VGND VPWR _10144_/S _10615_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout384 VGND VPWR fanout390/X _10347_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout362 VGND VPWR _10588_/S _10732_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout373 VGND VPWR _11162_/S _11170_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_74_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout395 VGND VPWR _10890_/A _11235_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_15620_ _15620_/Q clkload27/A _15620_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13196__313 VPWR VGND VPWR VGND _14471_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_12832_ VGND VPWR VPWR VGND _15565_/D _12831_/X _12830_/Y _12834_/C1 _10056_/Y _15565_/Q
+ sky130_fd_sc_hd__a32o_1
X_15551_ _15551_/Q clkload32/A _15551_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12763_ VGND VPWR VGND VPWR _15548_/D _10060_/A _15548_/Q _09976_/B _12762_/Y sky130_fd_sc_hd__o211a_1
XFILLER_43_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14502_ _14502_/Q _14502_/CLK _14502_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13237__354 VPWR VGND VPWR VGND _14512_/CLK clkload11/A sky130_fd_sc_hd__inv_2
X_15482_ _15482_/Q _15482_/CLK _15482_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11714_ VPWR VGND VPWR VGND _11713_/X _12473_/A _12491_/B1 _11714_/X sky130_fd_sc_hd__a21o_1
X_12694_ VGND VPWR VPWR VGND _12695_/B _12693_/Y _12694_/S _12685_/Y sky130_fd_sc_hd__mux2_1
X_14433_ hold987/A _14433_/CLK _14433_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11645_ VGND VPWR VPWR VGND _11645_/X hold414/A _11964_/S hold200/A sky130_fd_sc_hd__mux2_1
X_11576_ VGND VPWR VPWR VGND _11580_/B hold611/A _12086_/S hold320/A sky130_fd_sc_hd__mux2_1
X_14364_ hold913/A _14364_/CLK _14364_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14295_ hold227/A _14295_/CLK _14295_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10527_ VGND VPWR VPWR VGND _10527_/X hold547/A _10627_/S hold472/A sky130_fd_sc_hd__mux2_1
XFILLER_13_1361 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10458_ VGND VPWR VGND VPWR _10458_/X _10486_/A1 _10454_/X _10457_/X _10704_/C1 sky130_fd_sc_hd__o211a_1
X_10389_ VGND VPWR VPWR VGND _10389_/X _14195_/Q _10390_/S hold252/A sky130_fd_sc_hd__mux2_1
X_12128_ VGND VPWR VGND VPWR _12128_/X _12156_/A1 _12124_/X _12127_/X _12202_/C1 sky130_fd_sc_hd__o211a_1
X_12059_ VGND VPWR VPWR VGND _12059_/X _14200_/Q _12219_/S hold181/A sky130_fd_sc_hd__mux2_1
XFILLER_77_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_53_706 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_80_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_761 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_463 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09270_ VGND VPWR VPWR VGND _14773_/D _09862_/A0 _09275_/S hold534/X sky130_fd_sc_hd__mux2_1
X_08221_ VPWR VGND VPWR VGND _07810_/A _15610_/Q _08249_/A2 _08230_/A _08218_/Y sky130_fd_sc_hd__a22o_1
X_08152_ VGND VPWR VPWR VGND _08152_/X _07563_/Y _08151_/Y _07596_/X _07591_/Y _07421_/A
+ sky130_fd_sc_hd__o2111a_1
X_07103_ VPWR VGND VPWR VGND _08880_/A _15152_/Q sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_9_clk clkload27/A clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_08083_ VGND VPWR _08083_/B _10063_/A _08083_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13902__1019 VPWR VGND VPWR VGND _15274_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_13030__147 VPWR VGND VPWR VGND _14273_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_08985_ VGND VPWR VGND VPWR hold945/A hold944/X _08985_/A2 _08984_/X _11337_/C1 sky130_fd_sc_hd__o211a_1
X_07936_ VPWR VGND VPWR VGND _15350_/Q _07560_/X _15139_/Q clone18/A _07936_/X sky130_fd_sc_hd__a22o_2
X_13678__795 VPWR VGND VPWR VGND _15018_/CLK clkload54/A sky130_fd_sc_hd__inv_2
XFILLER_29_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07867_ VPWR VGND VGND VPWR _07867_/A _07868_/B _07867_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_1298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_1359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07798_ VGND VPWR _07958_/D _07992_/B _07798_/A _07798_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_09606_ VGND VPWR VPWR VGND _14462_/D clone6/X _09619_/S hold378/X sky130_fd_sc_hd__mux2_1
X_09537_ VGND VPWR VPWR VGND _14525_/D fanout38/X _09537_/S hold311/X sky130_fd_sc_hd__mux2_1
X_09468_ VGND VPWR VPWR VGND _14588_/D fanout36/X _09478_/S hold237/X sky130_fd_sc_hd__mux2_1
XFILLER_11_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_24_496 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08419_ VGND VPWR _08418_/X _08735_/C _08419_/Y hold150/X VPWR VGND sky130_fd_sc_hd__o21ai_1
X_09399_ VGND VPWR VPWR VGND _14650_/D hold676/X _09406_/S fanout27/X sky130_fd_sc_hd__mux2_1
X_11430_ VGND VPWR VGND VPWR _11430_/X _14930_/Q _11303_/A _11431_/A2 sky130_fd_sc_hd__a21bo_1
X_11361_ VGND VPWR VPWR VGND _14852_/Q _11361_/X _14851_/Q sky130_fd_sc_hd__xor2_1
X_10312_ VGND VPWR VGND VPWR _10312_/X _11263_/C1 _10307_/X _10311_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_4_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11292_ VPWR VGND _14814_/D _11292_/B _11382_/S VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_65_1034 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10243_ VPWR VGND VGND VPWR _10243_/X _10911_/S _10243_/B sky130_fd_sc_hd__or2_1
X_10174_ VGND VPWR VPWR VGND _10174_/X _14349_/Q _10479_/S hold401/A sky130_fd_sc_hd__mux2_1
XFILLER_67_809 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout192 VGND VPWR _12684_/S _12581_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout170 VGND VPWR _12164_/A _12174_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_47_500 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout181 VGND VPWR _12721_/S _12396_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_14982_ hold457/A _14982_/CLK _14982_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_717 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_34_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12815_ VGND VPWR VGND VPWR _15561_/D _10056_/A _15561_/Q _07544_/B _12814_/X sky130_fd_sc_hd__o211a_1
X_15603_ _15603_/Q clkload32/A _15603_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15534_ _15534_/Q _15534_/CLK _15534_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12746_ VGND VPWR VGND VPWR _12746_/X _15512_/Q _12746_/A2 _11810_/S _12745_/X sky130_fd_sc_hd__o211a_1
X_13471__588 VPWR VGND VPWR VGND _14746_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_15465_ VGND VPWR VGND VPWR _15465_/Q _15465_/D clkload53/A sky130_fd_sc_hd__dfxtp_4
XFILLER_15_1401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12677_ VPWR VGND VGND VPWR _12658_/Y _12676_/X _12677_/A2 _15474_/Q _15474_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_15396_ _15396_/Q _15396_/CLK _15396_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_8_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14416_ hold816/A _14416_/CLK _14416_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11628_ VGND VPWR VPWR VGND _11628_/X _14863_/Q _11628_/S hold345/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14347_ hold851/A _14347_/CLK _14347_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11559_ VGND VPWR _11557_/B hold1288/X _11559_/Y _15439_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xhold607 hold607/X hold607/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 hold618/X hold618/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ _14278_/Q _14278_/CLK _14278_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14069__1186 VPWR VGND VPWR VGND _15488_/CLK clkload9/A sky130_fd_sc_hd__inv_2
Xhold629 hold629/X hold629/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_69_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13365__482 VPWR VGND VPWR VGND _14640_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
Xhold1307 hold1307/X _14845_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1318 hold1318/X _15587_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1329 hold1329/X _15586_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08770_ VGND VPWR VPWR VGND _15236_/D fanout6/X _08772_/S hold496/X sky130_fd_sc_hd__mux2_1
X_07721_ VPWR VGND VGND VPWR _15561_/Q _07938_/B _07721_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_555 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07652_ VPWR VGND VGND VPWR _07653_/B _07652_/A _07652_/B sky130_fd_sc_hd__or2_1
XFILLER_0_1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07583_ VGND VPWR VGND VPWR _07587_/B _09013_/B _08194_/B _10060_/C _08623_/B sky130_fd_sc_hd__o211ai_2
X_13712__829 VPWR VGND VPWR VGND _15052_/CLK clkload45/A sky130_fd_sc_hd__inv_2
XFILLER_0_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09322_ VGND VPWR VPWR VGND _14722_/D hold454/X _09327_/S clone54/X sky130_fd_sc_hd__mux2_1
XFILLER_34_794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_772 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09253_ VGND VPWR VPWR VGND _14790_/D _09272_/S fanout52/X hold1220/X sky130_fd_sc_hd__mux2_4
Xclone18 VGND VPWR clone18/X clone18/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_08204_ VPWR VGND VGND VPWR _15450_/Q _07369_/B _10074_/A1 _08204_/X sky130_fd_sc_hd__o21a_1
X_09184_ VGND VPWR VPWR VGND _14907_/D hold298/X _09188_/S fanout21/X sky130_fd_sc_hd__mux2_1
X_08135_ VPWR VGND _08136_/B _08135_/B _08135_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08066_ VPWR VGND VGND VPWR _08066_/A _08066_/B _08066_/Y sky130_fd_sc_hd__nor2_1
X_13606__723 VPWR VGND VPWR VGND _14946_/CLK clkload11/A sky130_fd_sc_hd__inv_2
XFILLER_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08968_ VGND VPWR VPWR VGND _08969_/B _07549_/A _09906_/A hold791/A sky130_fd_sc_hd__mux2_1
X_14188__906 _14188_/D _14188__906/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08899_ VGND VPWR VGND VPWR _15143_/D hold1364/X _08902_/B _08898_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
X_07919_ VPWR VGND VPWR VGND _08007_/A _07982_/B _07385_/Y _07942_/C sky130_fd_sc_hd__a21oi_1
X_10930_ VGND VPWR VGND VPWR _10930_/X _10927_/X _10929_/X _11235_/A1 _10930_/C1 sky130_fd_sc_hd__a211o_1
X_10861_ VGND VPWR VPWR VGND _10861_/X _14496_/Q _10885_/S hold405/A sky130_fd_sc_hd__mux2_1
X_12600_ VGND VPWR VGND VPWR _12600_/X _12599_/X _12598_/X _12375_/S _12863_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_73_1336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10792_ VGND VPWR VGND VPWR _10792_/X _10791_/X _10790_/X _11205_/A _11217_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_73_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12531_ VGND VPWR VPWR VGND _12531_/X _14501_/Q _12539_/S hold470/A sky130_fd_sc_hd__mux2_1
XFILLER_9_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15250_ _15250_/Q _15250_/CLK _15250_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12462_ VGND VPWR VPWR VGND _12462_/X _12459_/X _12476_/S _12458_/X sky130_fd_sc_hd__mux2_1
X_11413_ VPWR VGND VPWR VGND _11410_/Y _14857_/Q _14858_/Q _11413_/X sky130_fd_sc_hd__a21o_1
X_14201_ _14201_/Q _14201_/CLK _14201_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15181_ hold726/A _15181_/CLK _15181_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12393_ VGND VPWR VPWR VGND _12393_/X _14465_/Q _12408_/S _14753_/Q sky130_fd_sc_hd__mux2_1
X_11344_ VGND VPWR VGND VPWR _11344_/X _11421_/B _11343_/Y _11316_/Y _11327_/A sky130_fd_sc_hd__o211a_1
X_13349__466 VPWR VGND VPWR VGND _14624_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_14132_ hold239/A _14132_/CLK _14132_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11275_ VPWR VGND VGND VPWR _11557_/B _15438_/Q _11555_/B sky130_fd_sc_hd__or2_1
XFILLER_4_654 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_1364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_10_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10226_ VGND VPWR VGND VPWR _10226_/X _15002_/Q _11003_/A2 _10225_/X _10985_/S sky130_fd_sc_hd__o211a_1
XFILLER_80_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10157_ VGND VPWR VPWR VGND _10157_/X hold882/A _10169_/B hold333/A sky130_fd_sc_hd__mux2_1
XFILLER_0_860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14965_ hold932/A _14965_/CLK _14965_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10088_ VGND VPWR VGND VPWR _10088_/X _10614_/A1 _10084_/X _10087_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
X_14896_ hold649/A _14896_/CLK _14896_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13901__1018 VPWR VGND VPWR VGND _15273_/CLK clkload14/A sky130_fd_sc_hd__inv_2
X_12729_ VGND VPWR VPWR VGND _12729_/X _12726_/X _12735_/S _12725_/X sky130_fd_sc_hd__mux2_1
X_15517_ hold511/A _15517_/CLK _15517_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15448_ _15448_/Q clkload37/A _15448_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_50_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15379_ hold712/A _15379_/CLK _15379_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold426 hold426/X hold426/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 hold415/X hold415/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 hold404/X hold404/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ VGND VPWR VPWR VGND _14131_/D _09956_/S _09940_/S _09937_/Y sky130_fd_sc_hd__mux2_1
X_12964__81 VPWR VGND VPWR VGND _14207_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
Xhold459 hold459/X hold459/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 hold437/X hold437/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 hold448/X hold448/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09871_ VPWR VGND VGND VPWR hold212/X _09871_/Y _09888_/S sky130_fd_sc_hd__nand2_1
Xhold1104 hold1104/X _14528_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 hold1115/X _15131_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08822_ VGND VPWR VPWR VGND _15191_/D fanout77/X _08846_/S hold537/X sky130_fd_sc_hd__mux2_1
Xhold1148 _11549_/A _15435_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 _15104_/D _09000_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 hold1137/X _15337_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ VGND VPWR VPWR VGND _15253_/D fanout69/X _08776_/S hold893/X sky130_fd_sc_hd__mux2_1
XFILLER_6_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1159 _11551_/A _15436_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07704_ VGND VPWR VPWR VGND _07706_/B _15592_/Q _07807_/S _07519_/B sky130_fd_sc_hd__mux2_1
X_13142__259 VPWR VGND VPWR VGND _14417_/CLK clkload54/A sky130_fd_sc_hd__inv_2
XFILLER_39_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_864 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_2_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08684_ VGND VPWR VPWR VGND _08684_/X _14397_/Q _08684_/S _14381_/Q sky130_fd_sc_hd__mux2_1
XFILLER_38_374 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07635_ VPWR VGND VPWR VGND _07634_/Y _07619_/B _07984_/S _07635_/X sky130_fd_sc_hd__a21o_1
X_07566_ VGND VPWR VGND VPWR _07480_/Y _08687_/S _07566_/B sky130_fd_sc_hd__nand2b_2
XFILLER_41_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09305_ VGND VPWR VPWR VGND _14736_/D _09862_/A0 _09310_/S hold390/X sky130_fd_sc_hd__mux2_1
X_09236_ VPWR VGND VPWR VGND _14806_/Q hold280/X hold1305/X _09237_/C sky130_fd_sc_hd__a21oi_1
X_07497_ _08566_/B _07492_/A _07496_/Y _07492_/B _07456_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_13036__153 VPWR VGND VPWR VGND _14279_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09167_ VGND VPWR VPWR VGND _14924_/D hold329/X _09191_/S fanout86/X sky130_fd_sc_hd__mux2_1
XFILLER_79_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_79_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08118_ _10063_/C _11899_/A _07358_/B _08116_/A _08081_/A _08117_/X VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__o311a_1
X_09098_ VGND VPWR VPWR VGND _14997_/D hold359/X _09124_/S fanout83/X sky130_fd_sc_hd__mux2_1
X_13840__957 VPWR VGND VPWR VGND _15212_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_08049_ VPWR VGND VPWR VGND _08293_/A3 _07271_/B _08048_/X _08049_/Y sky130_fd_sc_hd__a21oi_1
Xhold971 hold971/X hold971/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold960 hold960/X hold960/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 hold982/X hold982/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ VPWR VGND VPWR VGND _11059_/X _11181_/A1 _11058_/X _11060_/Y sky130_fd_sc_hd__a21oi_1
X_10011_ VPWR VGND VPWR VGND _10010_/C _15619_/Q hold1301/X _10012_/B sky130_fd_sc_hd__a21oi_1
Xhold993 hold993/X hold993/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13693__810 VPWR VGND VPWR VGND _15033_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_62_1037 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14750_ hold620/A _14750_/CLK _14750_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_45_812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13734__851 VPWR VGND VPWR VGND _15106_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_11962_ VGND VPWR VPWR VGND _11966_/B hold794/A _11964_/S hold788/A sky130_fd_sc_hd__mux2_1
XFILLER_28_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14068__1185 VPWR VGND VPWR VGND _15487_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_11893_ VPWR VGND VGND VPWR _11894_/S _11889_/X _12189_/C1 _11893_/X sky130_fd_sc_hd__o21a_1
X_10913_ VGND VPWR VPWR VGND _10914_/B _10912_/Y _10987_/S _10904_/Y sky130_fd_sc_hd__mux2_1
X_14681_ hold440/A _14681_/CLK _14681_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10844_ VGND VPWR VPWR VGND _10844_/X hold846/A _10850_/S hold786/A sky130_fd_sc_hd__mux2_1
X_15302_ _15302_/Q _15302_/CLK _15302_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10775_ VGND VPWR VPWR VGND _10775_/X hold726/A _10850_/S hold432/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12514_ VPWR VGND VGND VPWR _12514_/X hold386/A _12671_/S sky130_fd_sc_hd__or2_1
XFILLER_51_1442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_768 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15233_ hold279/A _15233_/CLK _15233_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12445_ VGND VPWR VPWR VGND _12445_/X hold772/A _12623_/S hold346/A sky130_fd_sc_hd__mux2_1
X_12376_ VPWR VGND VPWR VGND _12375_/X _12373_/X _12374_/X _12376_/X _12376_/B2 sky130_fd_sc_hd__a22o_1
X_15164_ hold498/A _15164_/CLK _15164_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11327_ VGND VPWR _14827_/D _11327_/B _11327_/A _11327_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_15095_ _15095_/Q clkload36/A _15095_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11258_ VGND VPWR VGND VPWR _11258_/X _15512_/Q _11262_/A2 _11257_/X _10851_/A sky130_fd_sc_hd__o211a_1
X_10209_ VPWR VGND VPWR VGND _10208_/X _11237_/A1 _10207_/X _10209_/Y sky130_fd_sc_hd__a21oi_1
X_11189_ VGND VPWR VGND VPWR _11189_/X _11186_/X _11188_/X _11189_/A1 _11245_/A1 sky130_fd_sc_hd__a211o_1
X_13477__594 VPWR VGND VPWR VGND _14752_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_14948_ hold894/A _14948_/CLK _14948_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14879_ _14879_/Q _14879_/CLK _14879_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07420_ VPWR VGND _07421_/A _07420_/X _08286_/B VPWR VGND sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07351_ VPWR VGND VPWR VGND _07351_/Y _07899_/B sky130_fd_sc_hd__inv_2
XFILLER_17_1348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07282_ VPWR VGND _07288_/A _07285_/B _15463_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_09021_ VPWR VGND VGND VPWR _15479_/Q _15477_/Q _08935_/A _09022_/B sky130_fd_sc_hd__o21a_1
Xhold201 hold201/X hold201/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/X hold212/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/X hold234/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/X hold223/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold278/X hold278/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold256 hold256/X hold256/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/X hold267/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/X hold245/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ VPWR VGND VPWR VGND _14136_/Q _09923_/D _14135_/Q _14140_/Q _09931_/C sky130_fd_sc_hd__or4_1
Xfanout703 VPWR VGND _08448_/B _08425_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout714 VGND VPWR _11490_/S _11475_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xhold289 hold289/X hold289/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout725 VGND VPWR _11974_/A1 _12602_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout747 VGND VPWR _07572_/X _08232_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout758 VPWR VGND _08604_/B2 _07524_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout736 VGND VPWR _09975_/Y _12834_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09854_ VGND VPWR VPWR VGND _14168_/D hold820/X _09864_/S fanout20/X sky130_fd_sc_hd__mux2_1
Xfanout769 VGND VPWR _07420_/X _07881_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_08805_ VGND VPWR VPWR VGND _15204_/D fanout6/X _08806_/S hold303/X sky130_fd_sc_hd__mux2_1
X_13718__835 VPWR VGND VPWR VGND _15058_/CLK clkload48/A sky130_fd_sc_hd__inv_2
XFILLER_27_801 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09785_ VGND VPWR VPWR VGND _14264_/D fanout19/X _09790_/S hold383/X sky130_fd_sc_hd__mux2_1
X_08736_ VGND VPWR _08738_/B _14766_/Q _09938_/C _14763_/Q VPWR VGND sky130_fd_sc_hd__o21ai_2
XANTENNA_107 fanout424/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08667_ VGND VPWR VGND VPWR _08667_/X _08667_/A2 _08700_/B1 _15291_/Q _08666_/X sky130_fd_sc_hd__a211o_1
XANTENNA_118 _12694_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07618_ VPWR VGND VPWR VGND _07908_/B1 _15635_/Q _07952_/A2 _07629_/A _15599_/Q sky130_fd_sc_hd__a22o_1
XFILLER_74_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08598_ VGND VPWR _08598_/B _08598_/Y _08598_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_70_1317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07549_ VPWR VGND VGND VPWR _07549_/A _07549_/B _07556_/B sky130_fd_sc_hd__nor2_1
X_10560_ VPWR VGND _10560_/X _10550_/X _10546_/X _10626_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
X_13270__387 VPWR VGND VPWR VGND _14545_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_09219_ VGND VPWR VPWR VGND _14874_/D hold1041/X _09231_/S fanout15/X sky130_fd_sc_hd__mux2_1
X_10491_ VGND VPWR VPWR VGND _10491_/X hold795/A _10521_/B hold651/A sky130_fd_sc_hd__mux2_1
X_12230_ VGND VPWR VGND VPWR _12230_/X _12227_/X _12229_/X _12230_/A1 _12230_/C1 sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_80_Right_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12161_ VGND VPWR VPWR VGND _12161_/X _14491_/Q _12183_/S hold683/A sky130_fd_sc_hd__mux2_1
X_13900__1017 VPWR VGND VPWR VGND _15272_/CLK clkload14/A sky130_fd_sc_hd__inv_2
X_11112_ VPWR VGND VGND VPWR _11112_/X _11112_/A _11112_/B sky130_fd_sc_hd__or2_1
Xhold790 hold790/X hold790/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12092_ VGND VPWR VPWR VGND _12092_/X _12089_/X _12100_/S _12088_/X sky130_fd_sc_hd__mux2_1
X_11043_ VPWR VGND VPWR VGND _11042_/X _11247_/A _12713_/B1 _11043_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_476 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13164__281 VPWR VGND VPWR VGND _14439_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_14802_ _14802_/Q clkload46/A _14802_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_58_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14733_ hold297/A _14733_/CLK _14733_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11945_ VGND VPWR VGND VPWR _11945_/X _11944_/X _11943_/X _11948_/S _12189_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_44_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14664_ _14664_/Q _14664_/CLK _14664_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11876_ VPWR VGND VGND VPWR _11876_/X hold169/A _11876_/B sky130_fd_sc_hd__or2_1
X_10827_ VGND VPWR VGND VPWR _10827_/X hold829/A _11215_/A2 _10826_/X _11086_/C1 sky130_fd_sc_hd__o211a_1
X_13511__628 VPWR VGND VPWR VGND _14786_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_14595_ hold269/A _14595_/CLK _14595_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10758_ VGND VPWR VPWR VGND _10758_/X hold908/A _10835_/B hold183/A sky130_fd_sc_hd__mux2_1
XFILLER_41_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_594 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15216_ _15216_/Q _15216_/CLK _15216_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10689_ VGND VPWR VGND VPWR _10689_/X _10686_/X _10688_/X _10698_/A1 _10693_/B1 sky130_fd_sc_hd__a211o_1
X_12428_ VGND VPWR VPWR VGND _12428_/X hold552/A _12651_/S hold339/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1256 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12359_ VGND VPWR VGND VPWR _12359_/X _12356_/X _12358_/X _12375_/S _12376_/B2 sky130_fd_sc_hd__a211o_1
X_15147_ _15147_/Q _15147_/CLK _15147_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12934__51 VPWR VGND VPWR VGND _14177_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_15078_ _15078_/Q clkload16/A _15078_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13405__522 VPWR VGND VPWR VGND _14680_/CLK clkload18/A sky130_fd_sc_hd__inv_2
XFILLER_68_712 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09570_ VGND VPWR VPWR VGND _14495_/D hold847/X _09587_/S fanout46/X sky130_fd_sc_hd__mux2_1
XFILLER_27_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08521_ VPWR VGND VGND VPWR _08553_/A2 hold923/X _08503_/Y _15324_/Q hold924/A _11398_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08452_ VPWR VGND VGND VPWR _08452_/X _15350_/Q _08488_/B sky130_fd_sc_hd__or2_1
XFILLER_63_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07403_ VPWR VGND VGND VPWR _07403_/X _07403_/A _07665_/C sky130_fd_sc_hd__or2_1
XFILLER_24_848 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08383_ VGND VPWR VPWR VGND _15394_/D fanout77/X _08405_/S hold930/X sky130_fd_sc_hd__mux2_1
XFILLER_17_1101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07334_ _07410_/B _07153_/B _15475_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_07265_ VPWR VGND VGND VPWR _14393_/Q _07230_/S _07265_/B1 _07267_/B sky130_fd_sc_hd__o21a_1
X_09004_ VPWR VGND VGND VPWR _09007_/A _09004_/B _09004_/Y sky130_fd_sc_hd__nor2_1
X_07196_ VPWR VGND VGND VPWR _08083_/A _07196_/B _07197_/A sky130_fd_sc_hd__nor2_1
X_14067__1184 VPWR VGND VPWR VGND _15486_/CLK clkload11/A sky130_fd_sc_hd__inv_2
X_09906_ VPWR VGND VGND VPWR _09906_/A _09906_/Y _09906_/B sky130_fd_sc_hd__nand2_1
Xfanout533 VGND VPWR _12282_/S _12689_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout500 VGND VPWR _12149_/S _12043_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout511 VGND VPWR _12409_/B _12408_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout522 VGND VPWR _12446_/B _12651_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13148__265 VPWR VGND VPWR VGND _14423_/CLK clkload10/A sky130_fd_sc_hd__inv_2
Xfanout544 VPWR VGND VGND VPWR _08034_/B1 clone18/A sky130_fd_sc_hd__buf_12
Xfanout566 _09449_/S _09441_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout555 VPWR VGND _09825_/S _09799_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout577 _09376_/S _09346_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout599 _08811_/S _08780_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout588 VPWR VGND _09055_/S _09056_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_09837_ VGND VPWR VPWR VGND _14185_/D hold594/X _09861_/S clone133/X sky130_fd_sc_hd__mux2_1
X_09768_ VGND VPWR VPWR VGND _14281_/D fanout85/X _09795_/S hold557/X sky130_fd_sc_hd__mux2_1
X_08719_ VGND VPWR VGND VPWR _15274_/D hold915/X _08721_/A2 _08718_/X _11294_/A sky130_fd_sc_hd__o211a_1
XFILLER_70_921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11730_ VGND VPWR VPWR VGND _11730_/X _11727_/X _12396_/S _11726_/X sky130_fd_sc_hd__mux2_1
X_09699_ VGND VPWR VPWR VGND _09710_/S fanout81/X hold1227/X _14344_/D sky130_fd_sc_hd__mux2_2
XFILLER_42_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11661_ VGND VPWR VPWR VGND _11661_/X _14349_/Q _11965_/S hold401/A sky130_fd_sc_hd__mux2_1
XFILLER_30_807 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14380_ VGND VPWR VGND VPWR _14380_/Q _14380_/D clkload7/A sky130_fd_sc_hd__dfxtp_4
X_11592_ VGND VPWR VGND VPWR _11592_/X _11591_/X _11590_/X _11625_/S _12099_/C1 sky130_fd_sc_hd__a211o_1
X_10612_ VGND VPWR VPWR VGND _10612_/X _14457_/Q _10612_/S _14745_/Q sky130_fd_sc_hd__mux2_1
XFILLER_23_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10543_ VGND VPWR VPWR VGND _10543_/X hold887/A _10554_/S hold504/A sky130_fd_sc_hd__mux2_1
X_13846__963 VPWR VGND VPWR VGND _15218_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_15001_ _15001_/Q _15001_/CLK _15001_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10474_ VPWR VGND VGND VPWR _10474_/X hold356/A _10484_/B sky130_fd_sc_hd__or2_1
XFILLER_29_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12213_ VGND VPWR VPWR VGND _12214_/B _12212_/Y _12213_/S _12204_/Y sky130_fd_sc_hd__mux2_1
X_12144_ VGND VPWR VGND VPWR _12144_/X _12143_/X _12142_/X _12156_/A1 _12202_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_2_752 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12075_ VGND VPWR VPWR VGND _12075_/X hold372/A _12227_/S hold701/A sky130_fd_sc_hd__mux2_1
XFILLER_65_715 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11026_ VPWR VGND VGND VPWR _11026_/X hold371/A _11175_/S sky130_fd_sc_hd__or2_1
XFILLER_80_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15696_ VPWR VGND uo_out[1] _15696_/A VPWR VGND sky130_fd_sc_hd__buf_2
X_14716_ hold418/A _14716_/CLK _14716_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11928_ VPWR VGND VGND VPWR _11928_/X hold158/A _12043_/B sky130_fd_sc_hd__or2_1
X_11859_ VGND VPWR VPWR VGND _11859_/X hold486/A _12117_/B hold447/A sky130_fd_sc_hd__mux2_1
X_14647_ hold472/A _14647_/CLK _14647_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_18 _09660_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_14578_ hold173/A _14578_/CLK _14578_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_29 _14408_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_18_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_53_1389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_70_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_64_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07952_ VPWR VGND VPWR VGND _15624_/Q _07952_/A2 _07953_/C _08002_/B1 _15588_/Q _07951_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07883_ VPWR VGND VPWR VGND _07882_/X _07881_/Y _07883_/B1 _07890_/B sky130_fd_sc_hd__a21oi_1
X_09622_ VGND VPWR VPWR VGND _14446_/D _09622_/A1 _09622_/S hold937/X sky130_fd_sc_hd__mux2_1
X_09553_ VGND VPWR VPWR VGND _14509_/D _09691_/A0 _09553_/S hold188/X sky130_fd_sc_hd__mux2_1
X_13789__906 VPWR VGND VPWR VGND _15161_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08504_ VPWR VGND VGND VPWR _14766_/Q _09912_/A _08508_/A sky130_fd_sc_hd__nor2_1
X_09484_ VGND VPWR VPWR VGND _14572_/D fanout99/X _09485_/S hold342/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13533__650 VPWR VGND VPWR VGND _14864_/CLK clkload23/A sky130_fd_sc_hd__inv_2
X_08435_ VGND VPWR VGND VPWR _15359_/D hold1236/X _08458_/B _08434_/X _11382_/S sky130_fd_sc_hd__o211a_1
XFILLER_51_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08366_ VGND VPWR VPWR VGND _15407_/D hold612/X _08366_/S fanout5/X sky130_fd_sc_hd__mux2_1
X_07317_ VPWR VGND VPWR VGND _07694_/A _07693_/B sky130_fd_sc_hd__inv_2
XFILLER_32_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08297_ VPWR VGND VPWR VGND _08174_/Y _14835_/Q _08296_/X _08297_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07248_ VGND VPWR VPWR VGND _08117_/A _08135_/B _08135_/A _07248_/A _07249_/B sky130_fd_sc_hd__or4_4
X_07179_ VGND VPWR VGND VPWR _07182_/A _14396_/Q _07304_/A2 _07304_/B1 _15462_/Q sky130_fd_sc_hd__o211a_1
X_10190_ VPWR VGND _10190_/X _10180_/X _10176_/X _10626_/C1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
Xfanout341 VGND VPWR _11107_/S _10850_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout330 VPWR VGND _11186_/S _10964_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_13382__499 VPWR VGND VPWR VGND _14657_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
Xfanout374 VGND VPWR _11162_/S _11176_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout352 VPWR VGND _10144_/S _08195_/C VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout363 VPWR VGND _10588_/S _08195_/C VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout396 VGND VPWR fanout405/A _10890_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout385 VGND VPWR fanout390/X _10523_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_12831_ VPWR VGND VGND VPWR _12831_/X _12831_/A _12831_/B sky130_fd_sc_hd__or2_1
X_15550_ _15550_/Q clkload43/A _15550_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12762_ VGND VPWR _12788_/S _12761_/X _12762_/Y _08210_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_43_976 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12693_ VPWR VGND VPWR VGND _12692_/X _12703_/A1 _12691_/X _12693_/Y sky130_fd_sc_hd__a21oi_1
X_14501_ _14501_/Q _14501_/CLK _14501_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13276__393 VPWR VGND VPWR VGND _14551_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_15481_ hold956/A _15481_/CLK _15481_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11713_ VPWR VGND _11713_/X _11712_/X _11708_/X _12472_/S _11704_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14432_ hold823/A _14432_/CLK _14432_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11644_ VGND VPWR VPWR VGND _11644_/X hold957/A _11954_/S hold215/A sky130_fd_sc_hd__mux2_1
XFILLER_35_1020 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14363_ _14363_/Q _14363_/CLK _14363_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11575_ VPWR VGND VPWR VGND _11574_/X _12101_/A1 _11573_/X _11575_/Y sky130_fd_sc_hd__a21oi_1
X_14294_ hold410/A _14294_/CLK _14294_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10526_ VPWR VGND VGND VPWR _10507_/Y _10525_/X _10192_/B _14390_/Q _14390_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
X_10457_ VPWR VGND VGND VPWR _10457_/X _10467_/S _10457_/B sky130_fd_sc_hd__or2_1
XFILLER_6_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_48_1425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12904__21 VPWR VGND VPWR VGND _14146_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_10388_ VGND VPWR VPWR VGND _10388_/X hold951/A _10390_/S hold169/A sky130_fd_sc_hd__mux2_1
X_12127_ VPWR VGND VGND VPWR _12127_/X _12147_/S _12127_/B sky130_fd_sc_hd__or2_1
X_12058_ VGND VPWR VPWR VGND _12058_/X hold383/A _12219_/S hold514/A sky130_fd_sc_hd__mux2_1
X_11009_ VGND VPWR VPWR VGND _11009_/X hold900/A _11165_/S hold642/A sky130_fd_sc_hd__mux2_1
XFILLER_53_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_770 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13517__634 VPWR VGND VPWR VGND _14792_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
XFILLER_34_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14066__1183 VPWR VGND VPWR VGND _15485_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_08220_ VPWR VGND VPWR VGND _08220_/B _08220_/C _08220_/A _08220_/X sky130_fd_sc_hd__or3_1
X_08151_ VPWR VGND VGND VPWR _11440_/B _08151_/Y _08151_/B sky130_fd_sc_hd__nand2_1
X_07102_ VPWR VGND VPWR VGND _08458_/A _07102_/A sky130_fd_sc_hd__inv_2
X_08082_ VPWR VGND VPWR VGND _08102_/B _07196_/B _07355_/Y _08083_/B sky130_fd_sc_hd__a21oi_1
X_08984_ VGND VPWR VGND VPWR _08984_/X _08983_/A _08972_/A _15108_/Q _08983_/Y sky130_fd_sc_hd__a211o_1
XFILLER_69_873 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07935_ VPWR VGND VPWR VGND _15350_/Q _07560_/X _07935_/Y _15139_/Q clone19/X sky130_fd_sc_hd__a22oi_2
X_09605_ VGND VPWR VPWR VGND _14463_/D fanout47/X _09619_/S hold573/X sky130_fd_sc_hd__mux2_1
X_07866_ VPWR VGND VPWR VGND _15628_/Q _07952_/A2 _07870_/A _08002_/B1 _15592_/Q _07865_/Y
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07797_ VPWR VGND _07798_/C _07736_/B _07795_/C _15556_/Q _07733_/Y VGND VPWR sky130_fd_sc_hd__a31o_1
X_09536_ VGND VPWR VPWR VGND _14526_/D fanout41/X _09537_/S hold209/X sky130_fd_sc_hd__mux2_1
XFILLER_37_781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09467_ VGND VPWR VPWR VGND _14589_/D fanout40/X _09467_/S hold256/X sky130_fd_sc_hd__mux2_1
XFILLER_52_740 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08418_ VGND VPWR VGND VPWR _08418_/X _14808_/Q _14807_/Q _08413_/Y _08417_/Y sky130_fd_sc_hd__o211a_1
X_09398_ VGND VPWR VPWR VGND _14651_/D hold679/X _09414_/S fanout31/X sky130_fd_sc_hd__mux2_1
XFILLER_36_1373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08349_ VGND VPWR VPWR VGND _15424_/D hold310/X _08356_/S fanout69/X sky130_fd_sc_hd__mux2_1
XFILLER_7_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11360_ VPWR VGND VPWR VGND _11398_/D _11368_/A sky130_fd_sc_hd__inv_2
X_13310__427 VPWR VGND VPWR VGND _14585_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_10311_ VGND VPWR VGND VPWR _10311_/X _10310_/X _10309_/X _10315_/S _11259_/C1 sky130_fd_sc_hd__a211o_1
X_11291_ VGND VPWR VPWR VGND _11292_/B _14814_/Q _11299_/S _14382_/Q sky130_fd_sc_hd__mux2_1
X_10242_ VGND VPWR VPWR VGND _10242_/X hold693/A _10258_/B hold281/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10173_ VGND VPWR VPWR VGND _10173_/X hold896/A _10479_/S hold477/A sky130_fd_sc_hd__mux2_1
XFILLER_78_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout160 VPWR VGND _08933_/A _08932_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout171 VGND VPWR _12164_/A _11948_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout182 VPWR VGND _12721_/S _12367_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_14981_ hold331/A _14981_/CLK _14981_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13204__321 VPWR VGND VPWR VGND _14479_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
Xfanout193 VGND VPWR _12328_/S _12684_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_78_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15602_ _15602_/Q clkload19/A _15602_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12814_ VGND VPWR VGND VPWR _12814_/X _12812_/X _12813_/Y _12822_/A _09975_/A sky130_fd_sc_hd__a211o_1
X_15533_ hold305/A _15533_/CLK _15533_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12745_ VPWR VGND VGND VPWR _12745_/X _14538_/Q _12747_/S sky130_fd_sc_hd__or2_1
XFILLER_76_1197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15464_ VGND VPWR VGND VPWR _15464_/Q _15464_/D clkload54/A sky130_fd_sc_hd__dfxtp_4
X_12676_ VPWR VGND VPWR VGND _12675_/X _12658_/A _12713_/B1 _12676_/X sky130_fd_sc_hd__a21o_1
X_14415_ hold839/A _14415_/CLK _14415_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15395_ hold657/A _15395_/CLK _15395_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11627_ VGND VPWR VGND VPWR _11627_/X hold873/A _12040_/A2 _11638_/A1 _11626_/X sky130_fd_sc_hd__o211a_1
X_11558_ VPWR VGND VPWR VGND _11557_/Y _11277_/B _11341_/Y _15439_/D sky130_fd_sc_hd__a21oi_1
X_14346_ _14346_/Q _14346_/CLK _14346_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold608 hold608/X hold608/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ VGND VPWR VPWR VGND _10509_/X hold875/A _10516_/S hold870/A sky130_fd_sc_hd__mux2_1
Xhold619 hold619/X hold619/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ hold575/A _14277_/CLK _14277_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11489_ VGND VPWR VPWR VGND _15080_/D _11488_/X _11492_/S hold1424/X sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_891 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07720_ VPWR VGND VGND VPWR _07938_/A _15561_/Q _07721_/B sky130_fd_sc_hd__or2_1
Xhold1319 _10030_/A _15628_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1308 hold1308/X _15632_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_567 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07651_ VPWR VGND VGND VPWR _07665_/B _07665_/C _07665_/A _07652_/B sky130_fd_sc_hd__o21a_1
X_13751__868 VPWR VGND VPWR VGND _15123_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_07582_ VGND VPWR VPWR VGND _08623_/B _14153_/Q _08591_/B _10060_/C _08684_/S sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09321_ VGND VPWR VPWR VGND _14723_/D hold446/X _09342_/S fanout62/X sky130_fd_sc_hd__mux2_1
XFILLER_80_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_59_1395 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09252_ VGND VPWR VPWR VGND _14791_/D fanout57/X _09269_/S hold670/X sky130_fd_sc_hd__mux2_1
XFILLER_21_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclone19 VGND VPWR clone19/X clone20/X VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_08203_ VGND VPWR VGND VPWR _08203_/X _08240_/A _08202_/X _08200_/Y _08225_/C1 sky130_fd_sc_hd__o211a_1
X_09183_ VGND VPWR VPWR VGND _14908_/D hold430/X _09197_/S fanout26/X sky130_fd_sc_hd__mux2_1
X_08134_ VPWR VGND VPWR VGND _11440_/B _08295_/B _08134_/Y _07331_/A _08132_/A sky130_fd_sc_hd__a22oi_1
X_13645__762 VPWR VGND VPWR VGND _14985_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_08065_ VGND VPWR VGND VPWR _08065_/X _08277_/S _10062_/B _08063_/Y _08280_/B2 sky130_fd_sc_hd__o211a_1
XFILLER_27_1306 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_66_1399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12895__12 VPWR VGND VPWR VGND _14137_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_08967_ VGND VPWR VGND VPWR _15115_/D hold888/X _08985_/A2 _08966_/X _08943_/A sky130_fd_sc_hd__o211a_1
XFILLER_69_681 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08898_ VPWR VGND VGND VPWR _08898_/X _15143_/Q _08924_/B sky130_fd_sc_hd__or2_1
X_07918_ VGND VPWR _07918_/B _07918_/Y _07925_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_72_813 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07849_ VGND VPWR VPWR VGND _07849_/D _07849_/C _07849_/B _07849_/A clone55/A sky130_fd_sc_hd__or4_4
XFILLER_17_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10860_ VGND VPWR VPWR VGND _10860_/X _14624_/Q _11241_/S hold379/A sky130_fd_sc_hd__mux2_1
XFILLER_44_559 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09519_ VGND VPWR VPWR VGND _14540_/D fanout98/X _09520_/S hold647/X sky130_fd_sc_hd__mux2_1
X_10791_ VGND VPWR VPWR VGND _10791_/X hold490/A _10795_/S hold207/A sky130_fd_sc_hd__mux2_1
X_12530_ VGND VPWR VPWR VGND _12534_/B hold889/A _12652_/S hold365/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_49_Left_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_9_928 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12461_ VGND VPWR VGND VPWR _12461_/X _12489_/A1 _12457_/X _12460_/X _12485_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_12_467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11412_ VGND VPWR VGND VPWR _14857_/D _14857_/Q _11410_/Y _11411_/X _08541_/A sky130_fd_sc_hd__o211a_1
X_14200_ _14200_/Q _14200_/CLK _14200_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_12_489 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15180_ hold646/A _15180_/CLK _15180_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14131_ _14131_/Q _14131_/CLK _14131_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12392_ VGND VPWR VPWR VGND _12392_/X _14209_/Q _12408_/S _15217_/Q sky130_fd_sc_hd__mux2_1
X_11343_ VPWR VGND VPWR VGND _14822_/Q _11421_/D _11343_/Y _14833_/Q _11421_/A sky130_fd_sc_hd__a22oi_1
X_11274_ VPWR VGND VGND VPWR _11555_/B _15437_/Q _11274_/B sky130_fd_sc_hd__or2_1
X_10225_ VPWR VGND VGND VPWR _10225_/X hold406/A _11231_/S sky130_fd_sc_hd__or2_1
X_14065__1182 VPWR VGND VPWR VGND _15484_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_10156_ VPWR VGND VGND VPWR _10137_/Y _10155_/X _10710_/B _14380_/Q _14380_/D _11296_/A
+ sky130_fd_sc_hd__o221a_1
X_14212__930 _14212_/D _14212__930/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_47_320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10087_ VPWR VGND VGND VPWR _10087_/X _10613_/A _10087_/B sky130_fd_sc_hd__or2_1
X_14964_ hold813/A _14964_/CLK _14964_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14895_ hold483/A _14895_/CLK _14895_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_74_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13588__705 VPWR VGND VPWR VGND _14919_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_10989_ VPWR VGND VGND VPWR _10989_/X hold711/A _10994_/S sky130_fd_sc_hd__or2_1
X_12728_ VGND VPWR VGND VPWR _12728_/X _12737_/B1 _12724_/X _12727_/X _12739_/C1 sky130_fd_sc_hd__o211a_1
X_15516_ hold290/A _15516_/CLK _15516_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15447_ _15447_/Q clkload23/A _15447_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12659_ VPWR VGND VGND VPWR _12659_/X hold448/A _12661_/S sky130_fd_sc_hd__or2_1
X_13629__746 VPWR VGND VPWR VGND _14969_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_31_798 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_1243 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15378_ hold902/A _15378_/CLK _15378_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold405 hold405/X hold405/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 hold416/X hold416/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 hold427/X hold427/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ hold451/A _14329_/CLK _14329_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold438 hold438/X hold438/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 hold449/X hold449/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09870_ VPWR VGND VGND VPWR _09880_/B hold212/A _09888_/S sky130_fd_sc_hd__or2_1
XFILLER_48_1063 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08821_ VGND VPWR VPWR VGND _15192_/D fanout80/X _08846_/S hold510/X sky130_fd_sc_hd__mux2_1
Xhold1105 hold1105/X _15014_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ VGND VPWR VPWR VGND _15254_/D _08773_/S clone47/X hold1129/X sky130_fd_sc_hd__mux2_4
Xhold1127 hold1127/X _15290_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 hold1116/X _15279_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 hold1149/X _15249_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 hold1138/X _15209_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_802 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07703_ VPWR VGND VPWR VGND _07827_/B _07751_/C _12878_/A _07703_/A _07703_/X sky130_fd_sc_hd__or4_2
X_08683_ VGND VPWR VGND VPWR _15287_/D hold952/X _08701_/A2 _08682_/X _12085_/C1 sky130_fd_sc_hd__o211a_1
X_13181__298 VPWR VGND VPWR VGND _14456_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
XFILLER_66_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07634_ VPWR VGND VGND VPWR _07639_/A _07634_/Y _07634_/B sky130_fd_sc_hd__nand2_1
X_07565_ _08073_/B _07480_/Y _07566_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_34_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07496_ VPWR VGND VGND VPWR _07496_/A _08592_/B _07496_/Y _08586_/A sky130_fd_sc_hd__nand3_1
X_09304_ VGND VPWR VPWR VGND _14737_/D _09653_/A0 _09304_/S hold163/X sky130_fd_sc_hd__mux2_1
X_14089__1206 VPWR VGND VPWR VGND _15508_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_09235_ VPWR VGND VGND VPWR _09239_/B _09235_/B _14808_/D sky130_fd_sc_hd__nor2_1
X_13075__192 VPWR VGND VPWR VGND _14318_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_09166_ _14925_/D fanout91/X fanout87/X _09191_/S _09165_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09097_ _14998_/D fanout93/X fanout89/X _09122_/S _09096_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08117_ VPWR VGND VPWR VGND _08117_/B _08138_/A _08117_/A _08117_/X sky130_fd_sc_hd__or3_1
X_08048_ VPWR VGND VPWR VGND _07272_/D _08278_/B _08048_/X _08293_/B1 _15078_/Q _08047_/Y
+ sky130_fd_sc_hd__a221o_1
Xhold972 hold972/X hold972/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold950 hold950/X hold950/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 hold961/X hold961/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _15620_/Q _10014_/B _15619_/Q _10010_/C VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold994 hold994/X hold994/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 hold983/X hold983/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_415 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09999_ VPWR VGND _10003_/C _10000_/B _15615_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_49_629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13422__539 VPWR VGND VPWR VGND _14697_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_11961_ VPWR VGND VPWR VGND _11960_/X _12185_/A1 _11959_/X _11961_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_673 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13773__890 VPWR VGND VPWR VGND _15145_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_10912_ VPWR VGND VPWR VGND _10911_/X _11237_/A1 _10910_/X _10912_/Y sky130_fd_sc_hd__a21oi_1
X_11892_ VPWR VGND VGND VPWR _11892_/X _12180_/S _11892_/B sky130_fd_sc_hd__or2_1
X_14680_ hold799/A _14680_/CLK _14680_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10843_ VGND VPWR VPWR VGND _10843_/X hold817/A _10850_/S hold387/A sky130_fd_sc_hd__mux2_1
X_13316__433 VPWR VGND VPWR VGND _14591_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_10774_ VGND VPWR VGND VPWR _10774_/X _11218_/A1 _10769_/X _10773_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_44_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15301_ hold940/A _15301_/CLK _15301_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12513_ VGND VPWR VPWR VGND _12513_/X _12512_/X _12665_/S _12511_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15232_ hold221/A _15232_/CLK _15232_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12444_ VGND VPWR VGND VPWR _12444_/X _12656_/A1 _12439_/X _12443_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_12375_ VGND VPWR VPWR VGND _12375_/X _12372_/X _12375_/S _12371_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15163_ hold626/A _15163_/CLK _15163_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11326_ VPWR VGND VPWR VGND _11325_/Y _11313_/C _11317_/X _11327_/C sky130_fd_sc_hd__a21o_1
X_15094_ _15094_/Q clkload33/A _15094_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11257_ VPWR VGND VGND VPWR _11257_/X _14538_/Q _11261_/B sky130_fd_sc_hd__or2_1
XFILLER_80_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10208_ VGND VPWR VPWR VGND _10208_/X _10205_/X _10995_/S _10204_/X sky130_fd_sc_hd__mux2_1
X_11188_ VGND VPWR VGND VPWR _11188_/X _15028_/Q _11252_/A2 _11187_/X _11250_/S sky130_fd_sc_hd__o211a_1
X_10139_ VGND VPWR VGND VPWR _10139_/X _14863_/Q _10629_/A2 _10138_/X _10144_/S sky130_fd_sc_hd__o211a_1
X_14947_ hold637/A _14947_/CLK _14947_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14878_ _14878_/Q _14878_/CLK _14878_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_36_857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_63_698 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_1365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07350_ VPWR VGND VPWR VGND _07349_/X _07925_/A _07347_/X _07899_/B sky130_fd_sc_hd__a21o_1
X_13059__176 VPWR VGND VPWR VGND _14302_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_09020_ _09974_/A _15638_/Q _09024_/A _15479_/Q clone20/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_07281_ VPWR VGND VGND VPWR _14397_/Q _07304_/A2 _07304_/B1 _07285_/B sky130_fd_sc_hd__o21a_1
XFILLER_31_595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold202 hold202/X hold202/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/X hold235/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/X hold213/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/X hold224/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold257/X hold257/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 hold246/X hold246/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/X hold268/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout704 VPWR VGND _08458_/B _08425_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_09922_ VPWR VGND VGND VPWR hold1379/X _09919_/Y _09921_/Y _14136_/D sky130_fd_sc_hd__o21a_1
Xhold279 hold279/X hold279/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout715 VPWR VGND _11490_/S _10072_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout726 VPWR VGND _12491_/B1 _11974_/A1 VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout748 VGND VPWR _07563_/Y _10058_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout737 VGND VPWR _11458_/S _11476_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09853_ VGND VPWR VPWR VGND _14169_/D hold351/X _09867_/S fanout23/X sky130_fd_sc_hd__mux2_1
X_13757__874 VPWR VGND VPWR VGND _15129_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_08804_ VGND VPWR VPWR VGND _15205_/D fanout8/X _08814_/S hold478/X sky130_fd_sc_hd__mux2_1
Xfanout759 VGND VPWR _08002_/B1 _07908_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09784_ VGND VPWR VPWR VGND _14265_/D _09798_/S fanout23/X hold1215/X sky130_fd_sc_hd__mux2_4
X_08735_ _08734_/B _08851_/B _15262_/D _08735_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_13003__120 VPWR VGND VPWR VGND _14246_/CLK clkload53/A sky130_fd_sc_hd__inv_2
XANTENNA_119 _10893_/B1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_108 _10893_/B1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08666_ VPWR VGND VGND VPWR _08664_/X _08690_/S _08194_/Y _14403_/Q _08666_/X _08665_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_74_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08597_ VPWR VGND VGND VPWR _08597_/A _08598_/B _08597_/B sky130_fd_sc_hd__nand2_1
X_07617_ VGND VPWR VGND VPWR _07914_/B1 _07629_/B _07616_/X _07418_/B sky130_fd_sc_hd__o21ba_4
X_07548_ VGND VPWR VPWR VGND _07549_/B _07547_/Y _07523_/Y _07513_/X _07552_/B1 _15563_/Q
+ sky130_fd_sc_hd__a32o_1
XFILLER_14_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_74_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14064__1181 VPWR VGND VPWR VGND _15483_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_07479_ VGND VPWR VGND VPWR _07479_/Y _15446_/Q _07479_/A sky130_fd_sc_hd__xnor2_4
X_10490_ VGND VPWR VPWR VGND _10494_/B hold916/A _10520_/S hold632/A sky130_fd_sc_hd__mux2_1
X_09218_ VGND VPWR VPWR VGND _14875_/D hold1062/X _09229_/S fanout19/X sky130_fd_sc_hd__mux2_1
XFILLER_30_10 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09149_ VGND VPWR VPWR VGND _14949_/D fanout25/X _09163_/S hold801/X sky130_fd_sc_hd__mux2_1
X_12160_ VGND VPWR VPWR VGND _12164_/B hold639/A _12183_/S hold679/A sky130_fd_sc_hd__mux2_1
X_11111_ VGND VPWR VGND VPWR _11111_/X _11112_/A _11107_/X _11110_/X _11259_/C1 sky130_fd_sc_hd__o211a_1
Xhold791 hold791/X hold791/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold780 hold780/X hold780/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12091_ VGND VPWR VGND VPWR _12091_/X _12099_/A1 _12087_/X _12090_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
X_11042_ VPWR VGND _11042_/X _11041_/X _11037_/X _11246_/S _11033_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_7_1005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14801_ _14801_/Q clkload31/A _14801_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11944_ VGND VPWR VPWR VGND _11944_/X hold877/A _11964_/S hold497/A sky130_fd_sc_hd__mux2_1
X_14732_ hold309/A _14732_/CLK _14732_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11875_ VGND VPWR VPWR VGND _11875_/X hold811/A _11876_/B hold197/A sky130_fd_sc_hd__mux2_1
X_14663_ hold388/A _14663_/CLK _14663_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_17_356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10826_ VPWR VGND VGND VPWR _10826_/X hold317/A _10835_/B sky130_fd_sc_hd__or2_1
XFILLER_71_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13550__667 VPWR VGND VPWR VGND _14881_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_14594_ hold336/A _14594_/CLK _14594_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10757_ VGND VPWR VPWR VGND _10761_/B hold493/A _10835_/B hold505/A sky130_fd_sc_hd__mux2_1
X_10688_ VGND VPWR VGND VPWR _10688_/X hold943/A _10688_/A2 _10687_/X _10685_/S sky130_fd_sc_hd__o211a_1
X_15215_ hold274/A _15215_/CLK _15215_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12427_ VGND VPWR VPWR VGND _12431_/B hold670/A _12651_/S hold198/A sky130_fd_sc_hd__mux2_1
X_12358_ VGND VPWR VGND VPWR _12358_/X hold999/A _12861_/A1 _12373_/A _12357_/X sky130_fd_sc_hd__o211a_1
X_15146_ _15146_/Q _15146_/CLK _15146_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11309_ VGND VPWR VGND VPWR _14827_/Q _14825_/Q _14826_/Q _14828_/Q _11421_/A sky130_fd_sc_hd__and4bb_1
X_13444__561 VPWR VGND VPWR VGND _14719_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_12289_ VGND VPWR VPWR VGND _12289_/X _14430_/Q _12701_/S _14686_/Q sky130_fd_sc_hd__mux2_1
X_15077_ _15077_/Q clkload16/A _15077_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14088__1205 VPWR VGND VPWR VGND _15507_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_3_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08520_ VPWR VGND _15326_/D _08520_/B _11420_/S VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_48_492 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08451_ VGND VPWR VGND VPWR _15351_/D _15350_/Q _08448_/B _08450_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
X_12889__6 VPWR VGND VPWR VGND _14131_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_07402_ VGND VPWR _07173_/B _07681_/B _07665_/C _07086_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
X_08382_ VGND VPWR VPWR VGND _15395_/D fanout80/X _08405_/S hold657/X sky130_fd_sc_hd__mux2_1
X_07333_ VPWR VGND VGND VPWR _07574_/A _07333_/Y _10072_/A sky130_fd_sc_hd__nand2_4
X_07264_ VGND VPWR VGND VPWR _07262_/X _08010_/A _07264_/B sky130_fd_sc_hd__nand2b_2
X_09003_ VGND VPWR VGND VPWR _09003_/X hold1097/X _09015_/A2 _09002_/X _09017_/A sky130_fd_sc_hd__o211a_1
X_07195_ VPWR VGND VGND VPWR _07196_/B _07195_/A _08104_/A sky130_fd_sc_hd__or2_1
XFILLER_65_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09905_ VPWR VGND VPWR VGND _09904_/Y _08862_/C _09893_/A _09906_/B sky130_fd_sc_hd__a21o_1
Xfanout501 VGND VPWR _07568_/X _12149_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout523 VGND VPWR _12446_/B _12652_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout512 VPWR VGND _12409_/B _12726_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout545 VPWR VGND VGND VPWR clone20/A _08034_/B1 sky130_fd_sc_hd__buf_8
Xfanout556 _09827_/S _09830_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_59_735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout534 VGND VPWR fanout538/X _12282_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout589 VPWR VGND _09053_/S _09056_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_09836_ _14186_/D fanout94/X fanout90/X _09864_/S _09835_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xfanout578 _09275_/S _09268_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout567 VPWR VGND _09441_/S _09415_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_09767_ _14282_/D fanout91/X fanout87/X _09765_/Y _09766_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08718_ VPWR VGND VPWR VGND hold840/X _08523_/B _08718_/X _08728_/B1 _14385_/Q _08722_/C1
+ sky130_fd_sc_hd__a221o_1
X_09698_ VGND VPWR VPWR VGND _14345_/D fanout84/X _09725_/S hold513/X sky130_fd_sc_hd__mux2_1
X_08649_ VGND VPWR VGND VPWR _08714_/A2 _14382_/Q _08194_/B _08649_/X sky130_fd_sc_hd__o21ba_1
X_11660_ VGND VPWR VPWR VGND _11660_/X hold896/A _11965_/S hold477/A sky130_fd_sc_hd__mux2_1
X_11591_ VGND VPWR VPWR VGND _11591_/X hold860/A _12094_/S hold517/A sky130_fd_sc_hd__mux2_1
X_10611_ VGND VPWR VPWR VGND _10611_/X _14201_/Q _10612_/S _15209_/Q sky130_fd_sc_hd__mux2_1
XFILLER_23_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13387__504 VPWR VGND VPWR VGND _14662_/CLK clkload52/A sky130_fd_sc_hd__inv_2
X_10542_ VGND VPWR VGND VPWR _10542_/X _10704_/C1 _10537_/X _10541_/X _10469_/S sky130_fd_sc_hd__o211a_1
XFILLER_41_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_41_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_565 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10473_ VGND VPWR VPWR VGND _10473_/X _10472_/X _10677_/S _10471_/X sky130_fd_sc_hd__mux2_1
X_15000_ _15000_/Q _15000_/CLK _15000_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12212_ VPWR VGND VPWR VGND _12211_/X _12212_/A1 _12210_/X _12212_/Y sky130_fd_sc_hd__a21oi_1
X_13428__545 VPWR VGND VPWR VGND _14703_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_12143_ VGND VPWR VPWR VGND _12143_/X hold828/A _12155_/S hold576/A sky130_fd_sc_hd__mux2_1
X_12074_ VGND VPWR VGND VPWR _12074_/X _12230_/C1 _12069_/X _12073_/X _12222_/C1 sky130_fd_sc_hd__o211a_1
X_11025_ VPWR VGND VGND VPWR _11247_/A _11025_/B _11025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_1239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_66_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14715_ hold409/A _14715_/CLK _14715_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15695_ VPWR VGND uo_out[0] _15695_/A VPWR VGND sky130_fd_sc_hd__buf_4
X_12995__112 VPWR VGND VPWR VGND _14238_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_11927_ VGND VPWR VPWR VGND _11927_/X hold765/A _12043_/B hold191/A sky130_fd_sc_hd__mux2_1
X_11858_ VGND VPWR VGND VPWR _11858_/X _15488_/Q _12188_/A2 _12106_/S _11857_/X sky130_fd_sc_hd__o211a_1
X_14646_ hold632/A _14646_/CLK _14646_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14577_ hold349/A _14577_/CLK _14577_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10809_ VPWR VGND VPWR VGND _10806_/X _11215_/C1 _10808_/X _10809_/X sky130_fd_sc_hd__a21o_1
XANTENNA_19 _09834_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_11789_ VPWR VGND VGND VPWR _11770_/Y _11788_/X _10192_/B _15450_/Q _15450_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
X_15129_ _15129_/Q _15129_/CLK _15129_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07951_ VPWR VGND VPWR VGND _07950_/Y _07810_/A _07939_/Y _07951_/X _12833_/A sky130_fd_sc_hd__a22o_1
XFILLER_64_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14063__1180 VPWR VGND VPWR VGND _15482_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_07882_ VPWR VGND VGND VPWR _07333_/Y _10075_/A _07876_/A _07879_/X _07882_/X sky130_fd_sc_hd__o22a_1
X_13221__338 VPWR VGND VPWR VGND _14496_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_09621_ VGND VPWR VPWR VGND _14447_/D _09829_/A1 _09622_/S hold693/X sky130_fd_sc_hd__mux2_1
XFILLER_7_1380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09552_ VGND VPWR VPWR VGND _14510_/D _09690_/A0 _09552_/S hold275/X sky130_fd_sc_hd__mux2_1
X_08503_ VPWR VGND VPWR VGND _08503_/Y _08503_/A sky130_fd_sc_hd__inv_2
XFILLER_23_1194 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09483_ VGND VPWR VPWR VGND _14573_/D _09726_/A1 _09485_/S hold200/X sky130_fd_sc_hd__mux2_1
X_08434_ VPWR VGND VGND VPWR _08434_/X _15359_/Q _08486_/B sky130_fd_sc_hd__or2_1
X_13869__986 VPWR VGND VPWR VGND _15241_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_23_145 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_71_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08365_ VGND VPWR VPWR VGND _15408_/D hold699/X _08366_/S fanout10/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07316_ VPWR VGND VPWR VGND _07693_/B _07316_/A _07316_/B sky130_fd_sc_hd__or2_2
X_08296_ VPWR VGND VPWR VGND _15153_/Q clone20/X _08296_/X _07560_/X _15332_/Q _08173_/Y
+ sky130_fd_sc_hd__a221o_1
X_13115__232 VPWR VGND VPWR VGND _14358_/CLK clkload11/A sky130_fd_sc_hd__inv_2
X_07247_ VGND VPWR VGND VPWR _07195_/A _07190_/B _07197_/A _07243_/X _07249_/A _07188_/X
+ sky130_fd_sc_hd__a221oi_2
X_07178_ VGND VPWR _07304_/A2 _07304_/B1 _07180_/B _14396_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xfanout320 VGND VPWR _10924_/B _10919_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout331 VGND VPWR _11068_/S _11179_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_21_Left_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout342 VGND VPWR fanout349/X _11107_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout364 VPWR VGND _08195_/C fanout382/X VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout375 VPWR VGND _11162_/S fanout381/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout353 VGND VPWR _10288_/S _10510_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout386 VGND VPWR fanout390/X _10634_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09819_ VGND VPWR VPWR VGND _14233_/D fanout23/X _09833_/S hold184/X sky130_fd_sc_hd__mux2_1
Xfanout397 VGND VPWR _11252_/C1 _11189_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_12830_ VPWR VGND VGND VPWR _12831_/A _12830_/Y _12830_/B sky130_fd_sc_hd__nand2_1
X_13813__930 VPWR VGND VPWR VGND _15185_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_12761_ VPWR VGND VGND VPWR _08208_/X _10079_/X _08200_/B _12789_/A _12761_/X _10060_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15480_ _15480_/Q _15480_/CLK _15480_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12692_ VGND VPWR VPWR VGND _12692_/X _12689_/X _12698_/S _12688_/X sky130_fd_sc_hd__mux2_1
X_14500_ hold900/A _14500_/CLK _14500_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11712_ VGND VPWR VGND VPWR _11712_/X _11709_/X _11711_/X _12489_/A1 _12722_/A1 sky130_fd_sc_hd__a211o_1
X_14431_ hold785/A _14431_/CLK _14431_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11643_ VGND VPWR VPWR VGND _11643_/X _14477_/Q _11954_/S hold636/A sky130_fd_sc_hd__mux2_1
XFILLER_30_627 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Left_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14087__1204 VPWR VGND VPWR VGND _15506_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_11574_ VGND VPWR VPWR VGND _11574_/X _11571_/X _12098_/A _11570_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14362_ hold918/A _14362_/CLK _14362_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14293_ hold176/A _14293_/CLK _14293_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10525_ VPWR VGND VPWR VGND _10524_/X _10507_/A _12047_/B1 _10525_/X sky130_fd_sc_hd__a21o_1
X_10456_ VGND VPWR VPWR VGND _10456_/X hold877/A _10464_/S hold497/A sky130_fd_sc_hd__mux2_1
X_13662__779 VPWR VGND VPWR VGND _15002_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_10387_ VGND VPWR VPWR VGND _10391_/B hold811/A _10390_/S hold197/A sky130_fd_sc_hd__mux2_1
X_12126_ VGND VPWR VPWR VGND _12126_/X hold745/A _12149_/S hold218/A sky130_fd_sc_hd__mux2_1
X_12057_ VGND VPWR VPWR VGND _12061_/B hold574/A _12219_/S hold302/A sky130_fd_sc_hd__mux2_1
X_11008_ VGND VPWR VPWR VGND _11012_/B hold579/A _11175_/S hold592/A sky130_fd_sc_hd__mux2_1
X_13556__673 VPWR VGND VPWR VGND _14887_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XFILLER_46_782 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_1389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_741 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_443 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13972__1089 VPWR VGND VPWR VGND _15344_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_14629_ hold889/A _14629_/CLK _14629_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08150_ VGND VPWR VPWR VGND _15521_/D _09685_/A0 _08267_/S hold271/X sky130_fd_sc_hd__mux2_1
XFILLER_21_649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07101_ VPWR VGND VPWR VGND _08448_/A _07101_/A sky130_fd_sc_hd__inv_2
X_08081_ VPWR VGND VGND VPWR _08081_/A _08102_/B _08081_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08983_ VPWR VGND VGND VPWR _08983_/A _08983_/B _08983_/Y sky130_fd_sc_hd__nor2_1
X_07934_ VGND VPWR VPWR VGND _15532_/D fanout41/X _07954_/S hold261/X sky130_fd_sc_hd__mux2_1
X_07865_ VPWR VGND VGND VPWR _07886_/A _07865_/B _07865_/Y sky130_fd_sc_hd__nor2_1
X_09604_ VGND VPWR VPWR VGND _09622_/S fanout48/X hold1232/X _14464_/D sky130_fd_sc_hd__mux2_2
X_07796_ VGND VPWR VPWR VGND _07958_/C _08037_/A _08056_/B _07795_/X _08057_/A _07738_/X
+ sky130_fd_sc_hd__o2111a_1
X_09535_ VGND VPWR VPWR VGND _14527_/D fanout44/X _09549_/S hold228/X sky130_fd_sc_hd__mux2_1
X_09466_ VGND VPWR VPWR VGND _14590_/D clone44/A _09467_/S hold207/X sky130_fd_sc_hd__mux2_1
XFILLER_25_977 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08417_ VPWR VGND VGND VPWR _14807_/Q _08415_/Y _08416_/Y _14808_/Q _08417_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_52_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09397_ VGND VPWR VPWR VGND _14652_/D hold319/X _09406_/S fanout36/X sky130_fd_sc_hd__mux2_1
X_08348_ VGND VPWR VPWR VGND _15425_/D _08372_/S hold1156/X fanout73/X sky130_fd_sc_hd__mux2_4
XFILLER_71_1254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_32_1238 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_32_1227 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08279_ VPWR VGND VPWR VGND _08293_/A3 _15066_/Q _08293_/B1 _08279_/X _07226_/Y sky130_fd_sc_hd__a22o_1
X_10310_ VGND VPWR VPWR VGND _10310_/X _14545_/Q _11098_/S hold349/A sky130_fd_sc_hd__mux2_1
X_11290_ VPWR VGND _14813_/D _11290_/B _11290_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_10241_ VGND VPWR VPWR VGND _10241_/X _14191_/Q _10919_/S hold264/A sky130_fd_sc_hd__mux2_1
X_10172_ VGND VPWR VGND VPWR _10172_/X _10704_/C1 _10167_/X _10171_/X _10469_/S sky130_fd_sc_hd__o211a_1
X_13499__616 VPWR VGND VPWR VGND _14774_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_14980_ hold335/A _14980_/CLK _14980_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout161 VPWR VGND _11542_/A _11341_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout150 VGND VPWR _08507_/X _08686_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout172 VPWR VGND _12164_/A _12180_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout183 VPWR VGND _12367_/S _12373_/A VPWR VGND sky130_fd_sc_hd__buf_4
X_13243__360 VPWR VGND VPWR VGND _14518_/CLK clkload11/A sky130_fd_sc_hd__inv_2
XFILLER_74_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout194 VGND VPWR _12373_/A _12328_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_15601_ _15601_/Q clkload32/A _15601_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12813_ VPWR VGND VGND VPWR _12822_/A _12813_/B _12813_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15532_ hold261/A _15532_/CLK _15532_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12744_ VGND VPWR VGND VPWR _12744_/X _12741_/X _12743_/X _12748_/A1 _12744_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_42_273 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15463_ _15463_/Q clkload53/A _15463_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_54_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12675_ VPWR VGND _12675_/X _12674_/X _12670_/X _12731_/S _12666_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15394_ hold930/A _15394_/CLK _15394_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14414_ hold833/A _14414_/CLK _14414_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11626_ VPWR VGND VGND VPWR _11626_/X hold483/A _11628_/S sky130_fd_sc_hd__or2_1
X_11557_ VPWR VGND VGND VPWR _11557_/A _11557_/Y _11557_/B sky130_fd_sc_hd__nand2_1
X_14345_ hold513/A _14345_/CLK _14345_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_8_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10508_ VGND VPWR VPWR VGND _10508_/X _14422_/Q _10516_/S hold815/A sky130_fd_sc_hd__mux2_1
Xhold609 hold609/X hold609/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ hold392/A _14276_/CLK _14276_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11488_ VGND VPWR VPWR VGND _11488_/X _11487_/X _11491_/S _15460_/Q sky130_fd_sc_hd__mux2_1
X_10439_ VPWR VGND VPWR VGND _10436_/X _10593_/A1 _10438_/X _10439_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12109_ VGND VPWR VPWR VGND _12109_/X _14876_/Q _12112_/S hold488/A sky130_fd_sc_hd__mux2_1
Xhold1309 hold1309/X _15617_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07650_ VPWR VGND VGND VPWR _07668_/A _07664_/A _07653_/A _07650_/X sky130_fd_sc_hd__o21a_1
X_07581_ VGND VPWR VPWR VGND _09013_/B _15545_/Q _08591_/B _10060_/C _07580_/Y sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13292__409 VPWR VGND VPWR VGND _14567_/CLK clkload42/A sky130_fd_sc_hd__inv_2
XFILLER_0_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09320_ VGND VPWR VPWR VGND _14724_/D hold561/X _09327_/S fanout65/X sky130_fd_sc_hd__mux2_1
X_09251_ VGND VPWR VPWR VGND _14792_/D fanout60/X _09272_/S hold661/X sky130_fd_sc_hd__mux2_1
XFILLER_22_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08202_ VGND VPWR VGND VPWR _08202_/X _08201_/A _08201_/B _08180_/C _08201_/Y sky130_fd_sc_hd__o211a_1
X_09182_ VGND VPWR VPWR VGND _14909_/D hold576/X _09188_/S fanout29/X sky130_fd_sc_hd__mux2_1
X_08133_ VGND VPWR VPWR VGND _08295_/B _08132_/A _08195_/A _10893_/B1 sky130_fd_sc_hd__mux2_1
X_08064_ VGND VPWR _08064_/B _10062_/B _08066_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13186__303 VPWR VGND VPWR VGND _14461_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
XFILLER_68_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13227__344 VPWR VGND VPWR VGND _14502_/CLK clkload52/A sky130_fd_sc_hd__inv_2
X_08966_ VPWR VGND VGND VPWR _08966_/X _08969_/A _08966_/B sky130_fd_sc_hd__or2_1
X_14086__1203 VPWR VGND VPWR VGND _15505_/CLK clkload37/A sky130_fd_sc_hd__inv_2
XFILLER_75_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08897_ VGND VPWR VGND VPWR _15144_/D _15143_/Q _08902_/B _08896_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
X_07917_ VPWR VGND VPWR VGND _07940_/B _07287_/Y _07288_/A _07918_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07848_ VPWR VGND VPWR VGND clone2/A _08286_/A clone17/X _07849_/D sky130_fd_sc_hd__a21oi_1
Xclone2 VGND VPWR clone2/X clone2/A VPWR VGND sky130_fd_sc_hd__clkbuf_1
X_09518_ VGND VPWR VPWR VGND _14541_/D _09726_/A1 _09520_/S hold414/X sky130_fd_sc_hd__mux2_1
X_07779_ VPWR VGND VPWR VGND _08187_/B _07756_/B _07754_/X _08153_/B sky130_fd_sc_hd__a21o_1
XFILLER_17_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_80_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10790_ VGND VPWR VGND VPWR _10790_/X _14334_/Q _11215_/A2 _10789_/X _11215_/C1 sky130_fd_sc_hd__o211a_1
X_09449_ VGND VPWR VPWR VGND _14603_/D fanout97/X _09449_/S hold876/X sky130_fd_sc_hd__mux2_1
XFILLER_33_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12460_ VPWR VGND VGND VPWR _12460_/X _12476_/S _12460_/B sky130_fd_sc_hd__or2_1
X_11411_ VGND VPWR VPWR VGND _11411_/X _14857_/Q _11410_/Y _11408_/A _11406_/C sky130_fd_sc_hd__o2bb2a_1
X_14042__1159 VPWR VGND VPWR VGND _15414_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_12391_ VGND VPWR VPWR VGND _12391_/X _14273_/Q _12408_/S _14305_/Q sky130_fd_sc_hd__mux2_1
X_11342_ VPWR VGND VGND VPWR _11342_/C _14827_/Q _14828_/Q _11421_/D sky130_fd_sc_hd__nor3_1
X_14130_ _14130_/Q _14130_/CLK _14130_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11273_ VPWR VGND VGND VPWR _11274_/B _11273_/A _11551_/B sky130_fd_sc_hd__or2_1
X_10224_ VGND VPWR VPWR VGND _10224_/X hold842/A _11231_/S hold614/A sky130_fd_sc_hd__mux2_1
XFILLER_4_689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10155_ VPWR VGND VPWR VGND _10154_/X _10618_/A _12121_/B1 _10155_/X sky130_fd_sc_hd__a21o_1
X_13971__1088 VPWR VGND VPWR VGND _15343_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_10086_ VGND VPWR VPWR VGND _10086_/X hold803/A _10271_/S hold199/A sky130_fd_sc_hd__mux2_1
X_14963_ _14963_/Q _14963_/CLK _14963_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_652 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_35_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14894_ hold369/A _14894_/CLK _14894_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_825 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13020__137 VPWR VGND VPWR VGND _14263_/CLK clkload14/A sky130_fd_sc_hd__inv_2
XFILLER_16_741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10988_ VPWR VGND VGND VPWR _11210_/A _10988_/B _10988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_774 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15515_ hold355/A _15515_/CLK _15515_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12727_ VPWR VGND VGND VPWR _12727_/X _12735_/S _12727_/B sky130_fd_sc_hd__or2_1
XFILLER_31_777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15446_ VGND VPWR VGND VPWR _15446_/Q _15446_/D clkload8/A sky130_fd_sc_hd__dfxtp_4
XFILLER_19_1380 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12658_ VPWR VGND VGND VPWR _12658_/A _12658_/B _12658_/Y sky130_fd_sc_hd__nor2_1
X_11609_ VPWR VGND VGND VPWR _11609_/X _12100_/S _11609_/B sky130_fd_sc_hd__or2_1
X_13668__785 VPWR VGND VPWR VGND _15008_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_12589_ VGND VPWR VPWR VGND _12589_/X _14438_/Q _12589_/S hold570/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_clk clkload19/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_15377_ hold802/A _15377_/CLK _15377_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold417 hold417/X hold417/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14328_ hold752/A _14328_/CLK _14328_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold406 hold406/X hold406/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14259_ hold951/A _14259_/CLK _14259_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold439 hold439/X hold439/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 hold428/X hold428/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08820_ VGND VPWR VPWR VGND _15193_/D fanout83/X _08844_/S hold841/X sky130_fd_sc_hd__mux2_1
Xhold1106 hold1106/X _14994_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 _11539_/A _15430_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 hold1128/X _14662_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1139 hold1139/X _14534_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_26_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08751_ VGND VPWR VPWR VGND _15255_/D fanout78/X _08773_/S hold348/X sky130_fd_sc_hd__mux2_1
X_07702_ VGND VPWR VGND VPWR _07810_/A _07807_/S _07827_/C _15572_/Q _07827_/A sky130_fd_sc_hd__and4_2
X_08682_ VPWR VGND VPWR VGND hold950/A _08562_/A _08682_/X _08691_/B1 _08681_/X _08688_/C1
+ sky130_fd_sc_hd__a221o_1
X_07633_ VPWR VGND VPWR VGND _07908_/B1 _15634_/Q _07952_/A2 _07643_/A _15598_/Q sky130_fd_sc_hd__a22o_1
XFILLER_54_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07564_ VPWR VGND VGND VPWR _07573_/A _07566_/B _07564_/B sky130_fd_sc_hd__nand2_1
X_07495_ VGND VPWR VPWR VGND _15454_/Q _08586_/A _15599_/Q sky130_fd_sc_hd__xor2_1
X_09303_ VGND VPWR VPWR VGND _14738_/D _09826_/A1 _09310_/S hold282/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1088 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09234_ VGND VPWR _09237_/B _09235_/B _09234_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_1322 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09165_ VPWR VGND VGND VPWR hold1360/X _09191_/S _09165_/Y sky130_fd_sc_hd__nand2b_1
X_08116_ VGND VPWR _08116_/B _08116_/Y _08116_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_14194__912 _14194_/D _14194__912/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_68_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09096_ VPWR VGND VGND VPWR hold1351/X _09124_/S _09096_/Y sky130_fd_sc_hd__nand2b_1
Xhold940 hold940/X hold940/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08047_ VPWR VGND VGND VPWR _08047_/A _08066_/B _08047_/Y sky130_fd_sc_hd__nor2_1
X_12955__72 VPWR VGND VPWR VGND _14198_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
Xhold973 hold973/X hold973/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 hold951/X hold951/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 hold962/X hold962/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold984 hold984/X hold984/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 hold995/X hold995/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09998_ VPWR VGND VGND VPWR _10000_/B _09998_/B _15614_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13461__578 VPWR VGND VPWR VGND _14736_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_08949_ VPWR VGND _15123_/D _08949_/B _11567_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_11960_ VGND VPWR VPWR VGND _11960_/X _11957_/X _12164_/A _11956_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_68_clk clkload12/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_10911_ VGND VPWR VPWR VGND _10911_/X _10908_/X _10911_/S _10907_/X sky130_fd_sc_hd__mux2_1
X_11891_ VGND VPWR VPWR VGND _11891_/X hold680/A _12191_/B hold271/A sky130_fd_sc_hd__mux2_1
X_10842_ VPWR VGND VPWR VGND _10839_/X _11086_/C1 _10841_/X _10842_/X sky130_fd_sc_hd__a21o_1
X_13355__472 VPWR VGND VPWR VGND _14630_/CLK clkload52/A sky130_fd_sc_hd__inv_2
X_10773_ VGND VPWR VGND VPWR _10773_/X _10772_/X _10771_/X _11092_/S _11217_/C1 sky130_fd_sc_hd__a211o_1
X_15300_ hold960/A _15300_/CLK _15300_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_40_541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12512_ VGND VPWR VPWR VGND _12512_/X hold955/A _12664_/S hold561/A sky130_fd_sc_hd__mux2_1
X_15231_ hold267/A _15231_/CLK _15231_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_60_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12443_ VGND VPWR VGND VPWR _12443_/X _12442_/X _12441_/X _12655_/S _12662_/C1 sky130_fd_sc_hd__a211o_1
X_15162_ _15162_/Q _15162_/CLK _15162_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_12374_ VPWR VGND VGND VPWR _12375_/S _12370_/X _12863_/A1 _12374_/X sky130_fd_sc_hd__o21a_1
X_11325_ VPWR VGND VGND VPWR _14827_/Q _14826_/Q _11325_/Y _14825_/Q sky130_fd_sc_hd__nand3_1
X_15093_ _15093_/Q clkload33/A _15093_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11256_ VGND VPWR VPWR VGND _11256_/X _15397_/Q _11261_/B _15544_/Q sky130_fd_sc_hd__mux2_1
XFILLER_5_987 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13702__819 VPWR VGND VPWR VGND _15042_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XFILLER_49_1395 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_45_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10207_ VGND VPWR VGND VPWR _10207_/X _11004_/A1 _10203_/X _10206_/X _11235_/C1 sky130_fd_sc_hd__o211a_1
X_11187_ VPWR VGND VGND VPWR _11187_/X hold340/A _11251_/B sky130_fd_sc_hd__or2_1
X_10138_ VPWR VGND VGND VPWR _10138_/X hold345/A _10140_/S sky130_fd_sc_hd__or2_1
X_10069_ VGND VPWR VPWR VGND _10069_/X _10066_/Y _07857_/B _07681_/Y _07622_/X _07621_/Y
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_leaf_59_clk clkload15/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_14946_ _14946_/Q _14946_/CLK _14946_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_47_195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14877_ _14877_/Q _14877_/CLK _14877_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1311 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07280_ VPWR VGND _07286_/B _07280_/B _15464_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_15429_ _15429_/Q _15429_/CLK _15429_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14085__1202 VPWR VGND VPWR VGND _15504_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_68_Left_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold225 hold225/X hold225/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 hold203/X hold203/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/X hold214/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ VPWR VGND VPWR VGND _09919_/Y _14136_/Q _09917_/A _09921_/Y sky130_fd_sc_hd__a21oi_1
Xhold258 hold258/X hold258/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold269/X hold269/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/X hold236/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/X hold247/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout705 VPWR VGND _08483_/A2 _08485_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout749 VGND VPWR _07534_/Y _08591_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout727 VPWR VGND _11974_/A1 _10053_/Y VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout738 VGND VPWR _11491_/S _11458_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout716 VGND VPWR _10072_/Y _11535_/C VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09852_ VGND VPWR VPWR VGND _14170_/D hold533/X _09865_/S fanout29/X sky130_fd_sc_hd__mux2_1
X_09783_ VGND VPWR VPWR VGND _14266_/D fanout27/X _09790_/S hold645/X sky130_fd_sc_hd__mux2_1
X_08803_ VGND VPWR VPWR VGND _15206_/D fanout13/X _08814_/S hold341/X sky130_fd_sc_hd__mux2_1
X_08734_ VGND VPWR _15263_/D _08734_/B _08735_/C _08851_/B VPWR VGND sky130_fd_sc_hd__and3_1
X_13298__415 VPWR VGND VPWR VGND _14573_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_14041__1158 VPWR VGND VPWR VGND _15413_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_6_1297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Left_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XANTENNA_109 _10737_/C1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_08665_ VPWR VGND VGND VPWR _14379_/Q _08194_/B _08728_/B1 _08665_/X sky130_fd_sc_hd__o21a_1
X_08596_ VGND VPWR VGND VPWR _15308_/D hold865/X _08628_/A2 _08595_/X _09000_/C1 sky130_fd_sc_hd__o211a_1
X_07616_ VPWR VGND VPWR VGND _15134_/Q _08034_/B1 hold728/A _07558_/B _07616_/X sky130_fd_sc_hd__a22o_2
XFILLER_42_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13339__456 VPWR VGND VPWR VGND _14614_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_07547_ VPWR VGND VGND VPWR _07547_/A _07547_/B _07547_/Y _07547_/C sky130_fd_sc_hd__nand3_1
XFILLER_35_1417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13970__1087 VPWR VGND VPWR VGND _15342_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_07478_ VPWR VGND VGND VPWR _07573_/A _15445_/Q _07571_/B sky130_fd_sc_hd__nand2_2
X_09217_ VGND VPWR VPWR VGND _14876_/D hold1067/X _09231_/S fanout26/X sky130_fd_sc_hd__mux2_1
X_09148_ VGND VPWR VPWR VGND _14950_/D fanout27/X _09161_/S hold828/X sky130_fd_sc_hd__mux2_1
X_09079_ VGND VPWR VPWR VGND _15014_/D hold1105/X _09092_/S fanout28/X sky130_fd_sc_hd__mux2_1
X_11110_ VPWR VGND VGND VPWR _11110_/X _11110_/A _11110_/B sky130_fd_sc_hd__or2_1
Xhold781 hold781/X hold781/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold770 hold770/X hold770/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12090_ VPWR VGND VGND VPWR _12090_/X _12098_/A _12090_/B sky130_fd_sc_hd__or2_1
XFILLER_77_703 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11041_ VGND VPWR VGND VPWR _11041_/X _11040_/X _11039_/X _11189_/A1 _11254_/C1 sky130_fd_sc_hd__a211o_1
Xhold792 hold792/X hold792/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14800_ _14800_/Q clkload47/A _14800_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11943_ VGND VPWR VGND VPWR _11943_/X hold717/A _12192_/A2 _11968_/S _11942_/X sky130_fd_sc_hd__o211a_1
X_14731_ hold165/A _14731_/CLK _14731_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_18_869 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14662_ _14662_/Q _14662_/CLK _14662_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11874_ VGND VPWR VPWR VGND _11874_/X _11873_/X _12174_/S _11872_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10825_ VGND VPWR VPWR VGND _10825_/X _10824_/X _11092_/S _10823_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_176 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13091__208 VPWR VGND VPWR VGND _14334_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_9_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14593_ _14593_/Q _14593_/CLK _14593_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10756_ VPWR VGND VPWR VGND _10755_/X _11218_/A1 _10754_/X _10756_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_872 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10687_ VPWR VGND VGND VPWR _10687_/X hold196/A _10687_/B sky130_fd_sc_hd__or2_1
X_15214_ hold172/A _15214_/CLK _15214_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12426_ VPWR VGND VPWR VGND _12425_/X _12656_/A1 _12424_/X _12426_/Y sky130_fd_sc_hd__a21oi_1
X_13132__249 VPWR VGND VPWR VGND _14375_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_15145_ _15145_/Q _15145_/CLK _15145_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12357_ VPWR VGND VGND VPWR _12357_/X _14304_/Q _12372_/S sky130_fd_sc_hd__or2_1
X_11308_ VGND VPWR VGND VPWR _14821_/D _14382_/Q _11303_/B _11307_/X _11308_/C1 sky130_fd_sc_hd__o211a_1
X_12288_ VPWR VGND VGND VPWR _12584_/A _12288_/B _12288_/Y sky130_fd_sc_hd__nor2_1
X_15076_ _15076_/Q clkload15/A _15076_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11239_ VGND VPWR VPWR VGND _11239_/X _14282_/Q _11251_/B _14314_/Q sky130_fd_sc_hd__mux2_1
XFILLER_23_1310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_23_1332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13026__143 VPWR VGND VPWR VGND _14269_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
XFILLER_3_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14929_ _14929_/Q clkload29/A _14929_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08450_ VPWR VGND VGND VPWR _08450_/X _15351_/Q _08488_/B sky130_fd_sc_hd__or2_1
X_13830__947 VPWR VGND VPWR VGND _15202_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_08381_ VGND VPWR VPWR VGND _15396_/D fanout83/X _08393_/S hold1021/X sky130_fd_sc_hd__mux2_1
X_07401_ VPWR VGND VGND VPWR _07679_/A _07681_/B _07401_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07332_ VPWR VGND VGND VPWR _15584_/Q _08198_/S _07332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13683__800 VPWR VGND VPWR VGND _15023_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_07263_ VPWR VGND VGND VPWR _07264_/B _15460_/Q _07263_/B sky130_fd_sc_hd__or2_1
X_09002_ VGND VPWR VGND VPWR _09002_/X _09007_/A _09016_/B1 _15102_/Q _09001_/Y sky130_fd_sc_hd__a211o_1
X_07194_ VPWR VGND VGND VPWR _07195_/A _08104_/A _08102_/A sky130_fd_sc_hd__nor2_1
X_13724__841 VPWR VGND VPWR VGND _15064_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_12925__42 VPWR VGND VPWR VGND _14168_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_09904_ VGND VPWR _09900_/A hold819/A _09904_/Y _14142_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
Xfanout524 VPWR VGND _12539_/S _12664_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout513 VGND VPWR fanout539/X _12726_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout502 VGND VPWR _12220_/S _12228_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout535 VGND VPWR _12577_/S _12578_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout546 VGND VPWR clone20/A _08252_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout557 _09830_/S _09799_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09835_ VPWR VGND VPWR VGND _09834_/B _09834_/A hold1430/X _09835_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_1337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout568 VPWR VGND _09443_/S _09446_/S VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout579 VPWR VGND _09268_/S _09241_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_09766_ VPWR VGND VGND VPWR _09766_/X _09766_/A _09792_/S sky130_fd_sc_hd__or2_1
X_08717_ VGND VPWR VGND VPWR _15275_/D hold895/X _08721_/A2 _08716_/X _08717_/C1 sky130_fd_sc_hd__o211a_1
X_09697_ _14346_/D fanout92/X fanout88/X _09695_/Y _09696_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
Xrebuffer40 VPWR VGND VPWR VGND rebuffer40/X rebuffer41/X sky130_fd_sc_hd__dlygate4sd1_1
X_08648_ VGND VPWR VGND VPWR _15296_/D hold907/X _08721_/A2 _08647_/X _11937_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_74_1252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_74_1241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08579_ VGND VPWR VGND VPWR _15311_/D hold1080/X _08628_/A2 _08578_/X _11337_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_1372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_1394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11590_ VGND VPWR VGND VPWR _11590_/X hold922/A _12040_/A2 _12099_/A1 _11589_/X sky130_fd_sc_hd__o211a_1
X_10610_ VGND VPWR VPWR VGND _10610_/X _14265_/Q _10612_/S hold170/A sky130_fd_sc_hd__mux2_1
X_10541_ VGND VPWR VGND VPWR _10541_/X _10538_/X _10540_/X _10705_/A _10706_/C1 sky130_fd_sc_hd__a211o_1
X_10472_ VGND VPWR VPWR VGND _10472_/X hold929/A _10472_/S hold572/A sky130_fd_sc_hd__mux2_1
X_12211_ VGND VPWR VPWR VGND _12211_/X _12208_/X _12221_/S _12207_/X sky130_fd_sc_hd__mux2_1
X_13467__584 VPWR VGND VPWR VGND _14742_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
XFILLER_29_1018 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12142_ VGND VPWR VGND VPWR _12142_/X _14877_/Q _12229_/A2 _12147_/S _12141_/X sky130_fd_sc_hd__o211a_1
X_12073_ VGND VPWR VGND VPWR _12073_/X _12072_/X _12071_/X _12221_/S _12226_/C1 sky130_fd_sc_hd__a211o_1
X_11024_ VGND VPWR VPWR VGND _11025_/B _11023_/Y _11246_/S _11015_/Y sky130_fd_sc_hd__mux2_1
XFILLER_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_739 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14084__1201 VPWR VGND VPWR VGND _15503_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_14714_ hold723/A _14714_/CLK _14714_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11926_ VGND VPWR VGND VPWR _11926_/X _12212_/A1 _11925_/X _11922_/X _12222_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_33_625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14645_ hold607/A _14645_/CLK _14645_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11857_ VPWR VGND VGND VPWR _11857_/X hold194/A _12117_/B sky130_fd_sc_hd__or2_1
XFILLER_60_477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10808_ VPWR VGND VPWR VGND _10807_/X _11213_/S _11217_/C1 _10808_/X sky130_fd_sc_hd__a21o_1
X_14576_ hold195/A _14576_/CLK _14576_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11788_ VPWR VGND VPWR VGND _11787_/X _12029_/A _12047_/B1 _11788_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_371 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10739_ VPWR VGND VGND VPWR _10739_/X hold316/A _10742_/S sky130_fd_sc_hd__or2_1
X_13708__825 VPWR VGND VPWR VGND _15048_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_14040__1157 VPWR VGND VPWR VGND _15412_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XFILLER_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12409_ VPWR VGND VGND VPWR _12409_/X hold168/A _12409_/B sky130_fd_sc_hd__or2_1
X_15128_ _15695_/A _15128_/CLK _15128_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07950_ VPWR VGND VPWR VGND _07950_/Y _07950_/A sky130_fd_sc_hd__inv_2
X_15059_ hold655/A _15059_/CLK _15059_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12891__8 VPWR VGND VPWR VGND _14133_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
XFILLER_64_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_60_1307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07881_ VPWR VGND VPWR VGND _07881_/A2 _15086_/Q _07880_/X _07881_/Y sky130_fd_sc_hd__a21oi_1
X_09620_ VGND VPWR VPWR VGND _14448_/D _09862_/A0 _09625_/S hold434/X sky130_fd_sc_hd__mux2_1
X_13260__377 VPWR VGND VPWR VGND _14535_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XFILLER_49_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_7_1392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09551_ VGND VPWR VPWR VGND _14511_/D _09689_/A0 _09552_/S hold167/X sky130_fd_sc_hd__mux2_1
XFILLER_23_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08502_ VPWR VGND _08502_/X _08502_/B _08507_/C VPWR VGND sky130_fd_sc_hd__and2_1
X_09482_ VGND VPWR VPWR VGND _14574_/D _09622_/A1 _09482_/S hold219/X sky130_fd_sc_hd__mux2_1
XFILLER_23_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08433_ VGND VPWR VGND VPWR _15360_/D hold1205/X _08458_/B _08432_/X _11388_/S sky130_fd_sc_hd__o211a_1
XFILLER_71_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08364_ VGND VPWR VPWR VGND _15409_/D hold650/X _08375_/S fanout14/X sky130_fd_sc_hd__mux2_1
XFILLER_32_691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07315_ VPWR VGND VGND VPWR _15469_/Q _07315_/B _07316_/B sky130_fd_sc_hd__nor2_1
X_13154__271 VPWR VGND VPWR VGND _14429_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_08295_ VPWR VGND VGND VPWR _08214_/A _08295_/B _08295_/Y sky130_fd_sc_hd__nand2b_1
X_07246_ VPWR VGND VPWR VGND _08116_/A _08136_/A _07243_/X _08100_/B sky130_fd_sc_hd__a21o_1
X_07177_ VGND VPWR VGND VPWR _07316_/A _07174_/Y _07663_/A _07314_/A sky130_fd_sc_hd__a21oi_2
XFILLER_30_1166 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13501__618 VPWR VGND VPWR VGND _14776_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
Xfanout321 VPWR VGND _10924_/B _11240_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout310 VGND VPWR _10735_/S _10743_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout332 VGND VPWR _11068_/S _11167_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout343 VGND VPWR _10795_/S _11204_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout354 VGND VPWR _10288_/S _10625_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout365 VGND VPWR _10985_/S _10995_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout387 VGND VPWR _10705_/A _10698_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout376 VGND VPWR fanout381/X _10851_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout398 VGND VPWR _11252_/C1 _11178_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09818_ VGND VPWR VPWR VGND _14234_/D fanout27/X _09825_/S hold159/X sky130_fd_sc_hd__mux2_1
XFILLER_28_920 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09749_ VGND VPWR VPWR VGND _14297_/D fanout23/X _09763_/S hold170/X sky130_fd_sc_hd__mux2_1
X_12760_ VPWR VGND VPWR VGND _12758_/Y _15547_/Q _12807_/B1 _15547_/D _12759_/X sky130_fd_sc_hd__a22o_1
X_12691_ VGND VPWR VGND VPWR _12691_/X _12256_/S _12687_/X _12690_/X _12702_/C1 sky130_fd_sc_hd__o211a_1
X_11711_ VGND VPWR VGND VPWR _11711_/X _15002_/Q _12488_/A2 _12470_/S _11710_/X sky130_fd_sc_hd__o211a_1
X_11642_ VGND VPWR VPWR VGND _11646_/B hold882/A _11950_/B hold333/A sky130_fd_sc_hd__mux2_1
X_14430_ _14430_/Q _14430_/CLK _14430_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14361_ hold949/A _14361_/CLK _14361_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11573_ VGND VPWR VGND VPWR _11573_/X _12099_/A1 _11569_/X _11572_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_11_897 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10524_ VPWR VGND _10524_/X _10523_/X _10519_/X _10469_/S _10515_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14292_ hold292/A _14292_/CLK _14292_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10455_ VGND VPWR VPWR VGND _10455_/X hold717/A _10464_/S hold177/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10386_ VPWR VGND VPWR VGND _10385_/X _10693_/B1 _10384_/X _10386_/Y sky130_fd_sc_hd__a21oi_1
X_12125_ VGND VPWR VPWR VGND _12125_/X hold700/A _12205_/S hold273/A sky130_fd_sc_hd__mux2_1
XFILLER_78_864 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_42_1004 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12056_ VPWR VGND VPWR VGND _12055_/X _12230_/C1 _12054_/X _12056_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11007_ VPWR VGND VGND VPWR _10988_/Y _11006_/X _12380_/B _14403_/Q _14403_/D _12492_/C1
+ sky130_fd_sc_hd__o221a_1
X_13097__214 VPWR VGND VPWR VGND _14340_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
XFILLER_0_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_55_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11909_ VGND VPWR VPWR VGND _11913_/B hold357/A _12227_/S hold338/A sky130_fd_sc_hd__mux2_1
X_13138__255 VPWR VGND VPWR VGND _14413_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_14628_ hold579/A _14628_/CLK _14628_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14559_ hold571/A _14559_/CLK _14559_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07100_ VGND VPWR VPWR VGND _08735_/C _07534_/A sky130_fd_sc_hd__clkinv_4
X_08080_ VGND VPWR _08080_/B _08080_/Y _08083_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_31_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13795__912 VPWR VGND VPWR VGND _15167_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_08982_ VGND VPWR VGND VPWR _15110_/D hold954/X _08985_/A2 _08981_/X _09017_/A sky130_fd_sc_hd__o211a_1
X_07933_ VGND VPWR VGND VPWR clone6/A _07932_/X _07933_/C _07933_/B _07933_/A sky130_fd_sc_hd__or4b_4
XFILLER_29_1371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07864_ VPWR VGND VGND VPWR _07865_/B _07864_/A _07864_/B sky130_fd_sc_hd__or2_1
X_13836__953 VPWR VGND VPWR VGND _15208_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_09603_ VGND VPWR VPWR VGND _14465_/D _09622_/S clone46/A hold1204/X sky130_fd_sc_hd__mux2_4
X_07795_ _07795_/X _07795_/C _07798_/A _07998_/B _07992_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_09534_ VGND VPWR VPWR VGND _09537_/S fanout49/X hold1104/X _14528_/D sky130_fd_sc_hd__mux2_2
X_09465_ VGND VPWR VPWR VGND _14591_/D fanout47/X _09467_/S hold526/X sky130_fd_sc_hd__mux2_1
XFILLER_52_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08416_ VPWR VGND VGND VPWR _14806_/Q hold280/X _08416_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_71_1233 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09396_ VGND VPWR VPWR VGND _14653_/D hold376/X _09408_/S fanout39/X sky130_fd_sc_hd__mux2_1
X_08347_ VGND VPWR VPWR VGND _15426_/D hold363/X _08356_/S clone146/X sky130_fd_sc_hd__mux2_1
X_08278_ VPWR VGND _08278_/X _08278_/B _08278_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_14083__1200 VPWR VGND VPWR VGND _15502_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_07229_ VPWR VGND _10061_/B _08278_/A _07229_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_10240_ VGND VPWR VPWR VGND _10240_/X hold703/A _10258_/B hold255/A sky130_fd_sc_hd__mux2_1
XFILLER_78_116 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10171_ VGND VPWR VGND VPWR _10171_/X _10168_/X _10170_/X _10486_/A1 _10693_/B1 sky130_fd_sc_hd__a211o_1
Xfanout140 VPWR VGND _08615_/B1 _08627_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout151 VPWR VGND _08503_/A _08502_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout173 VGND VPWR _08298_/A1 _12180_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout162 VGND VPWR _08522_/X _08728_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_74_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout195 VGND VPWR _07979_/X _12373_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13579__696 VPWR VGND VPWR VGND _14910_/CLK clkload21/A sky130_fd_sc_hd__inv_2
Xfanout184 VGND VPWR _12373_/A _12624_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_78_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15600_ _15600_/Q clkload44/A _15600_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12812_ VGND VPWR VPWR VGND _12812_/X _07950_/Y _12820_/B _07939_/Y sky130_fd_sc_hd__mux2_1
X_15531_ hold206/A _15531_/CLK _15531_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12743_ VGND VPWR VGND VPWR _12743_/X _15030_/Q _12743_/A2 _11810_/S _12742_/X sky130_fd_sc_hd__o211a_1
X_15462_ _15462_/Q clkload17/A _15462_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14413_ hold896/A _14413_/CLK _14413_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12674_ VGND VPWR VGND VPWR _12674_/X _12671_/X _12673_/X _12674_/A1 _12740_/A1 sky130_fd_sc_hd__a211o_1
X_15267__942 _15267_/D _15267__942/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_15393_ _15393_/Q _15393_/CLK _15393_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11625_ VGND VPWR VPWR VGND _11625_/X _11624_/X _11625_/S _11623_/X sky130_fd_sc_hd__mux2_1
X_11556_ VPWR VGND VPWR VGND _11555_/Y _11557_/B _11341_/Y _15438_/D sky130_fd_sc_hd__a21oi_1
XFILLER_7_610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14344_ _14344_/Q _14344_/CLK _14344_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14275_ hold507/A _14275_/CLK _14275_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10507_ VPWR VGND VGND VPWR _10507_/A _10507_/B _10507_/Y sky130_fd_sc_hd__nor2_1
X_11487_ VGND VPWR VPWR VGND _11487_/X _15081_/Q _11490_/S _15079_/Q sky130_fd_sc_hd__mux2_1
X_10438_ VPWR VGND VPWR VGND _10437_/X _10662_/S _10717_/C1 _10438_/X sky130_fd_sc_hd__a21o_1
X_13523__640 VPWR VGND VPWR VGND _14798_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_10369_ VPWR VGND VGND VPWR _10369_/X hold194/A _10632_/B sky130_fd_sc_hd__or2_1
XFILLER_61_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12108_ VGND VPWR VGND VPWR _12108_/X hold801/A _12188_/A2 _12119_/A1 _12107_/X sky130_fd_sc_hd__o211a_1
XFILLER_61_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12039_ VPWR VGND VGND VPWR _12039_/X hold546/A _12043_/B sky130_fd_sc_hd__or2_1
XFILLER_38_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07580_ VGND VPWR _07580_/B _07580_/Y _07580_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_53_528 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1226 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09250_ VGND VPWR VPWR VGND _14793_/D fanout65/X _09269_/S hold560/X sky130_fd_sc_hd__mux2_1
X_08201_ VPWR VGND VGND VPWR _08201_/A _08201_/B _08201_/Y _08201_/C sky130_fd_sc_hd__nand3_1
X_13372__489 VPWR VGND VPWR VGND _14647_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_09181_ VGND VPWR VPWR VGND _14910_/D hold337/X _09188_/S fanout33/X sky130_fd_sc_hd__mux2_1
X_08132_ VPWR VGND VPWR VGND _08132_/Y _08132_/A sky130_fd_sc_hd__inv_2
X_08063_ VPWR VGND VGND VPWR _08277_/S _08063_/Y _12790_/B sky130_fd_sc_hd__nand2_1
X_08965_ VGND VPWR VPWR VGND _08966_/B _07536_/X _09906_/A hold543/A sky130_fd_sc_hd__mux2_1
X_13266__383 VPWR VGND VPWR VGND _14541_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
XFILLER_57_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07916_ VPWR VGND VGND VPWR _07940_/B _07916_/A _07916_/B sky130_fd_sc_hd__or2_1
XFILLER_25_1021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08896_ VPWR VGND VGND VPWR _08896_/X _15144_/Q _08924_/B sky130_fd_sc_hd__or2_1
XFILLER_25_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13992__1109 VPWR VGND VPWR VGND _15364_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_07847_ VPWR VGND VPWR VGND _15629_/Q _07952_/A2 _07849_/C _07908_/B1 _15593_/Q _07846_/Y
+ sky130_fd_sc_hd__a221o_1
X_07778_ VPWR VGND VPWR VGND _08210_/B _08210_/A _07777_/A _08187_/B sky130_fd_sc_hd__a21o_1
X_09517_ VGND VPWR VPWR VGND _14542_/D _09622_/A1 _09517_/S hold503/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_80_892 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09448_ VGND VPWR VPWR VGND _14604_/D fanout98/X _09449_/S hold519/X sky130_fd_sc_hd__mux2_1
X_09379_ VGND VPWR VPWR VGND _14667_/D hold464/X _09379_/S fanout95/X sky130_fd_sc_hd__mux2_1
X_11410_ VPWR VGND VGND VPWR _11410_/A _11410_/B _11410_/Y sky130_fd_sc_hd__nor2_1
X_12390_ VGND VPWR VPWR VGND _12394_/B _14790_/Q _12408_/S _14241_/Q sky130_fd_sc_hd__mux2_1
X_11341_ VPWR VGND VGND VPWR _11341_/Y _11341_/A _11410_/A sky130_fd_sc_hd__nand2_2
X_11272_ VPWR VGND VGND VPWR _11551_/B _15435_/Q _11549_/B sky130_fd_sc_hd__or2_1
X_13507__624 VPWR VGND VPWR VGND _14782_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
XFILLER_4_679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10223_ VGND VPWR VGND VPWR _10223_/X _10220_/X _10222_/X _11004_/A1 _11235_/C1 sky130_fd_sc_hd__a211o_1
X_10154_ VPWR VGND _10154_/X _10153_/X _10149_/X _10617_/S _10145_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14962_ hold458/A _14962_/CLK _14962_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10085_ VGND VPWR VPWR VGND _10085_/X hold602/A _10271_/S hold160/A sky130_fd_sc_hd__mux2_1
XFILLER_78_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14893_ _14893_/Q _14893_/CLK _14893_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_71_870 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10987_ VGND VPWR VPWR VGND _10988_/B _10986_/Y _10987_/S _10978_/Y sky130_fd_sc_hd__mux2_1
XFILLER_16_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12726_ VGND VPWR VPWR VGND _12726_/X _14474_/Q _12726_/S _14762_/Q sky130_fd_sc_hd__mux2_1
X_15514_ hold233/A _15514_/CLK _15514_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15445_ VGND VPWR VGND VPWR _15445_/Q _15445_/D clkload6/A sky130_fd_sc_hd__dfxtp_4
X_12657_ VGND VPWR VPWR VGND _12658_/B _12656_/Y _12731_/S _12648_/Y sky130_fd_sc_hd__mux2_1
X_15376_ hold718/A _15376_/CLK _15376_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11608_ VGND VPWR VPWR VGND _11608_/X hold647/A _12097_/S hold342/A sky130_fd_sc_hd__mux2_1
X_12588_ VGND VPWR VGND VPWR _12588_/X _12587_/X _12586_/X _12588_/A1 _12748_/C1 sky130_fd_sc_hd__a211o_1
X_14327_ hold850/A _14327_/CLK _14327_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_11_1109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11539_ VPWR VGND VGND VPWR _11539_/A _11539_/Y _11539_/B sky130_fd_sc_hd__nand2_1
Xhold407 hold407/X hold407/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 hold418/X hold418/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ hold529/A _14258_/CLK _14258_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold429 hold429/X hold429/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14189_ _14189_/Q _14189_/CLK _14189_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1032 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13939__1056 VPWR VGND VPWR VGND _15311_/CLK clkload46/A sky130_fd_sc_hd__inv_2
XFILLER_39_801 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1129 hold1129/X _15254_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1107 hold1107/X _15013_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08750_ VGND VPWR VPWR VGND _15256_/D clone45/X _08773_/S hold247/X sky130_fd_sc_hd__mux2_1
Xhold1118 hold1118/X _14696_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08681_ VGND VPWR VPWR VGND _08681_/X _14398_/Q _08684_/S _14382_/Q sky130_fd_sc_hd__mux2_1
X_13300__417 VPWR VGND VPWR VGND _14575_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_07701_ VGND VPWR VPWR VGND _15537_/D fanout62/X _08251_/S hold204/X sky130_fd_sc_hd__mux2_1
X_07632_ VGND VPWR VGND VPWR clone17/X _07643_/B _07631_/X _07418_/B sky130_fd_sc_hd__o21ba_4
X_07563_ VPWR VGND VGND VPWR _07563_/A _07563_/B _07563_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09302_ VGND VPWR VPWR VGND _14739_/D _09825_/A1 _09302_/S hold615/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07494_ VPWR VGND _07494_/X _08592_/B _08592_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_21_211 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09233_ VGND VPWR _09237_/B hold280/A _14807_/Q _14806_/Q VPWR VGND sky130_fd_sc_hd__and3_1
X_09164_ VGND VPWR VPWR VGND _09198_/C _09198_/B _09486_/B _09164_/A _09164_/X sky130_fd_sc_hd__or4_4
XFILLER_33_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08115_ VPWR VGND VGND VPWR _08115_/A _08136_/A _08116_/B sky130_fd_sc_hd__nor2_1
X_09095_ VPWR VGND VPWR VGND _09095_/X _09729_/A _09095_/B sky130_fd_sc_hd__or2_2
X_08046_ VGND VPWR VGND VPWR _08046_/X _12794_/B _08045_/Y _08240_/A _07333_/Y sky130_fd_sc_hd__a211o_1
Xhold930 hold930/X hold930/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 hold963/X hold963/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 hold952/X hold952/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 hold941/X hold941/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/X hold985/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12970__87 VPWR VGND VPWR VGND _14213_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
Xhold996 hold996/X hold996/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 hold974/X hold974/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ VPWR VGND VPWR VGND _09996_/C _15613_/Q hold1342/X _09997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08948_ VPWR VGND VPWR VGND _08969_/A hold1439/X _08932_/X _08949_/B _15123_/Q sky130_fd_sc_hd__a22o_1
X_08879_ VGND VPWR VGND VPWR _15153_/D hold1387/X _08919_/A2 _08878_/X _11308_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_28_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_45_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10910_ VGND VPWR VGND VPWR _10910_/X _11189_/A1 _10906_/X _10909_/X _11254_/C1 sky130_fd_sc_hd__o211a_1
X_11890_ VGND VPWR VPWR VGND _11890_/X hold821/A _12191_/B hold381/A sky130_fd_sc_hd__mux2_1
X_10841_ VPWR VGND VPWR VGND _10840_/X _10315_/S _11096_/C1 _10841_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_870 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10772_ VGND VPWR VPWR VGND _10772_/X hold868/A _11091_/S hold452/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12511_ VGND VPWR VPWR VGND _12511_/X hold925/A _12664_/S hold469/A sky130_fd_sc_hd__mux2_1
X_15230_ hold484/A _15230_/CLK _15230_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12442_ VGND VPWR VPWR VGND _12442_/X _14885_/Q _12661_/S hold425/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15161_ hold151/A _15161_/CLK _15161_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12373_ VPWR VGND VGND VPWR _12373_/X _12373_/A _12373_/B sky130_fd_sc_hd__or2_1
X_11324_ VPWR VGND _11327_/B _11313_/C _14825_/Q _14826_/Q _14827_/Q VGND VPWR sky130_fd_sc_hd__a31o_1
X_15092_ _15092_/Q clkload33/A _15092_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_966 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13741__858 VPWR VGND VPWR VGND _15113_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_11255_ VGND VPWR VGND VPWR _11255_/X _11263_/C1 _11250_/X _11254_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
X_10206_ VPWR VGND VGND VPWR _10206_/X _10995_/S _10206_/B sky130_fd_sc_hd__or2_1
X_11186_ VGND VPWR VPWR VGND _11186_/X hold510/A _11186_/S hold624/A sky130_fd_sc_hd__mux2_1
X_13594__711 VPWR VGND VPWR VGND _14925_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_10137_ VPWR VGND VGND VPWR _10618_/A _10137_/B _10137_/Y sky130_fd_sc_hd__nor2_1
X_14945_ hold830/A _14945_/CLK _14945_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10068_ VGND VPWR VPWR VGND _10068_/X _10067_/X _07923_/B _07878_/X _07607_/Y _07410_/C
+ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_75_483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13635__752 VPWR VGND VPWR VGND _14975_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_39_1009 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14876_ _14876_/Q _14876_/CLK _14876_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_572 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12709_ VPWR VGND VGND VPWR _12709_/X hold359/A _12747_/S sky130_fd_sc_hd__or2_1
XFILLER_31_564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15428_ hold463/A _15428_/CLK _15428_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13991__1108 VPWR VGND VPWR VGND _15363_/CLK clkload32/A sky130_fd_sc_hd__inv_2
X_15359_ _15359_/Q _15359_/CLK _15359_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold226 hold226/X hold226/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/X hold215/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold204 hold204/X hold204/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ VGND VPWR VGND VPWR _09917_/A _09918_/X _09919_/Y _14137_/D sky130_fd_sc_hd__o21ba_1
Xhold248 hold248/X hold248/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold259/X hold259/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 hold237/X hold237/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout706 VGND VPWR _08425_/X _08485_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09851_ VGND VPWR VPWR VGND _14171_/D hold683/X _09867_/S fanout32/X sky130_fd_sc_hd__mux2_1
Xfanout739 VPWR VGND _11491_/S _09965_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout728 VGND VPWR _10192_/B _10710_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout717 VGND VPWR _10072_/Y _11529_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09782_ VGND VPWR VPWR VGND _14267_/D fanout31/X _09798_/S hold943/X sky130_fd_sc_hd__mux2_1
X_08802_ VGND VPWR VPWR VGND _15207_/D fanout16/X _08814_/S hold324/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08733_ VPWR VGND VGND VPWR _08733_/A _08853_/A _08851_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08664_ VPWR VGND VGND VPWR _08664_/X _14387_/Q _08664_/B sky130_fd_sc_hd__or2_1
X_08595_ VGND VPWR VGND VPWR _08595_/X _08617_/A _08615_/B1 _15307_/Q _08594_/Y sky130_fd_sc_hd__a211o_1
X_13378__495 VPWR VGND VPWR VGND _14653_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07615_ VGND VPWR VPWR VGND _15543_/D fanout83/X _07954_/S hold325/X sky130_fd_sc_hd__mux2_1
X_07546_ VPWR VGND VGND VPWR _07523_/B _07544_/X _07523_/Y _07545_/Y _07549_/A sky130_fd_sc_hd__o22a_1
XFILLER_35_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07477_ VGND VPWR VPWR VGND _07571_/B _15577_/Q _07477_/S _15590_/Q sky130_fd_sc_hd__mux2_1
XFILLER_50_895 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14202__920 _14202_/D _14202__920/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09216_ VGND VPWR VPWR VGND _14877_/D hold1102/X _09231_/S fanout28/X sky130_fd_sc_hd__mux2_1
XFILLER_10_737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09147_ VGND VPWR VPWR VGND _14951_/D fanout32/X _09163_/S hold992/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1205 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09078_ VGND VPWR VPWR VGND _15015_/D hold1049/X _09094_/S fanout34/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Left_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08029_ VPWR VGND VPWR VGND _15079_/Q _07420_/X _08029_/X _08293_/A3 _07268_/A _08028_/Y
+ sky130_fd_sc_hd__a221o_1
Xhold782 hold782/X hold782/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 hold771/X hold771/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_947 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold760 hold760/X hold760/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ VGND VPWR VPWR VGND _11040_/X hold627/A _11186_/S hold272/A sky130_fd_sc_hd__mux2_1
XFILLER_1_457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold793 hold793/X hold793/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14009__1126 VPWR VGND VPWR VGND _15381_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_79_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1460 hold1460/X hold923/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_612 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13619__736 VPWR VGND VPWR VGND _14959_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_79_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11942_ VPWR VGND VGND VPWR _11942_/X hold177/A _11950_/B sky130_fd_sc_hd__or2_1
XFILLER_45_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14730_ _14730_/Q _14730_/CLK _14730_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_17_325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11873_ VGND VPWR VPWR VGND _11873_/X hold569/A _11876_/B hold615/A sky130_fd_sc_hd__mux2_1
X_14661_ hold365/A _14661_/CLK _14661_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10824_ VGND VPWR VPWR VGND _10824_/X hold847/A _11093_/S hold767/A sky130_fd_sc_hd__mux2_1
X_14592_ hold254/A _14592_/CLK _14592_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13938__1055 VPWR VGND VPWR VGND _15310_/CLK clkload31/A sky130_fd_sc_hd__inv_2
XFILLER_38_1064 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10755_ VGND VPWR VPWR VGND _10755_/X _10752_/X _11205_/A _10751_/X sky130_fd_sc_hd__mux2_1
X_10686_ VGND VPWR VPWR VGND _10686_/X hold608/A _10687_/B hold185/A sky130_fd_sc_hd__mux2_1
X_15213_ hold277/A _15213_/CLK _15213_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13171__288 VPWR VGND VPWR VGND _14446_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_12425_ VGND VPWR VPWR VGND _12425_/X _12422_/X _12655_/S _12421_/X sky130_fd_sc_hd__mux2_1
X_12356_ VGND VPWR VPWR VGND _12356_/X _14789_/Q _12370_/S _14240_/Q sky130_fd_sc_hd__mux2_1
X_15144_ _15144_/Q _15144_/CLK _15144_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11307_ VPWR VGND VGND VPWR _11307_/X _14821_/Q _11307_/B sky130_fd_sc_hd__or2_1
X_12287_ VGND VPWR VPWR VGND _12288_/B _12286_/Y _12583_/S _12278_/Y sky130_fd_sc_hd__mux2_1
X_15075_ _15075_/Q clkload14/A _15075_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11238_ VGND VPWR VPWR VGND _11242_/B _14799_/Q _11251_/B _14250_/Q sky130_fd_sc_hd__mux2_1
X_11169_ VGND VPWR VGND VPWR _11169_/X _11178_/C1 _11165_/X _11168_/X _11180_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_49_962 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13065__182 VPWR VGND VPWR VGND _14308_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_14928_ _14928_/Q clkload29/A _14928_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14859_ _14859_/Q clkload26/A _14859_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08380_ _15397_/D fanout93/X fanout89/X _08378_/Y _08379_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07400_ _07401_/B _07315_/B _15469_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_1_1195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07331_ VPWR VGND VPWR VGND _08198_/S _07331_/A _08286_/B sky130_fd_sc_hd__or2_2
X_13412__529 VPWR VGND VPWR VGND _14687_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_07262_ VPWR VGND _07262_/X _07263_/B _15460_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_09001_ VPWR VGND VGND VPWR _09007_/A _09001_/B _09001_/Y sky130_fd_sc_hd__nor2_1
X_07193_ VPWR VGND VGND VPWR _15455_/Q _07355_/B _08104_/A sky130_fd_sc_hd__nor2_1
X_13763__880 VPWR VGND VPWR VGND _15135_/CLK clkload19/A sky130_fd_sc_hd__inv_2
X_09903_ VPWR VGND VPWR VGND _09902_/X _08860_/Y _09893_/Y _14142_/D hold1143/X sky130_fd_sc_hd__a22o_1
Xfanout514 VGND VPWR _12370_/S _12599_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout503 VGND VPWR _12220_/S _12219_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout536 VGND VPWR _12577_/S _12318_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout547 VPWR VGND clone20/A _07558_/Y VPWR VGND sky130_fd_sc_hd__buf_6
X_09834_ VPWR VGND VGND VPWR _09834_/Y _09834_/A _09834_/B sky130_fd_sc_hd__nand2_2
X_13306__423 VPWR VGND VPWR VGND _14581_/CLK clkload22/A sky130_fd_sc_hd__inv_2
Xfanout525 VGND VPWR _12446_/B _12664_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_12940__57 VPWR VGND VPWR VGND _14183_/CLK clkload42/A sky130_fd_sc_hd__inv_2
Xfanout569 _09446_/S _09415_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout558 _09728_/S _09721_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_55_921 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09765_ VPWR VGND VPWR VGND _09765_/Y _09792_/S sky130_fd_sc_hd__inv_2
Xrebuffer30 VPWR VGND VPWR VGND rebuffer30/X rebuffer31/X sky130_fd_sc_hd__dlygate4sd1_1
X_08716_ VPWR VGND VPWR VGND hold915/A _08523_/B _08716_/X _08728_/B1 _14386_/Q _08722_/C1
+ sky130_fd_sc_hd__a221o_1
X_09696_ VPWR VGND VGND VPWR _09696_/X _09696_/A _09725_/S sky130_fd_sc_hd__or2_1
Xrebuffer41 VPWR VGND VPWR VGND rebuffer41/X rebuffer42/X sky130_fd_sc_hd__dlygate4sd1_1
X_08647_ VPWR VGND VPWR VGND hold1450/X _08667_/A2 _08647_/X _08662_/B1 _08646_/X
+ _08700_/B1 sky130_fd_sc_hd__a221o_1
X_08578_ VGND VPWR VGND VPWR _08578_/X _08582_/A _08615_/B1 hold990/A _08577_/Y sky130_fd_sc_hd__a211o_1
XFILLER_74_1275 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07529_ VPWR VGND VPWR VGND _07551_/B _07551_/A _07433_/A _07545_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_1248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_50_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10540_ VGND VPWR VGND VPWR _10540_/X hold771/A _10583_/A2 _10539_/X _10703_/A sky130_fd_sc_hd__o211a_1
X_10471_ VGND VPWR VPWR VGND _10471_/X hold766/A _10484_/B hold849/A sky130_fd_sc_hd__mux2_1
X_12210_ VGND VPWR VGND VPWR _12210_/X _12230_/A1 _12206_/X _12209_/X _12226_/C1 sky130_fd_sc_hd__o211a_1
X_12141_ VPWR VGND VGND VPWR _12141_/X hold375/A _12205_/S sky130_fd_sc_hd__or2_1
Xhold590 hold590/X hold590/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12072_ VGND VPWR VPWR VGND _12072_/X _14875_/Q _12220_/S hold437/A sky130_fd_sc_hd__mux2_1
X_11023_ VPWR VGND VPWR VGND _11022_/X _11023_/A1 _11021_/X _11023_/Y sky130_fd_sc_hd__a21oi_1
X_13049__166 VPWR VGND VPWR VGND _14292_/CLK clkload16/A sky130_fd_sc_hd__inv_2
XFILLER_66_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1290 hold1290/X _15343_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13990__1107 VPWR VGND VPWR VGND _15362_/CLK clkload19/A sky130_fd_sc_hd__inv_2
XFILLER_46_976 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14713_ hold724/A _14713_/CLK _14713_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11925_ VGND VPWR VPWR VGND _11925_/X _11924_/X _11925_/S _11923_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_272 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11856_ VGND VPWR VGND VPWR _11856_/X _11853_/X _11855_/X _11958_/A _12175_/A1 sky130_fd_sc_hd__a211o_1
X_14644_ hold481/A _14644_/CLK _14644_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1337 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_53_1315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10807_ VGND VPWR VPWR VGND _10807_/X _14881_/Q _11216_/S _15417_/Q sky130_fd_sc_hd__mux2_1
X_14575_ hold461/A _14575_/CLK _14575_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11787_ VPWR VGND _11787_/X _11786_/X _11782_/X _12176_/S _11778_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10738_ VGND VPWR VPWR VGND _10738_/X hold633/A _10742_/S hold266/A sky130_fd_sc_hd__mux2_1
X_13747__864 VPWR VGND VPWR VGND _15119_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_10669_ VGND VPWR VGND VPWR _10669_/X hold936/A _10744_/A2 _10668_/X _10652_/S sky130_fd_sc_hd__o211a_1
X_12408_ VGND VPWR VPWR VGND _12408_/X hold610/A _12408_/S hold288/A sky130_fd_sc_hd__mux2_1
X_15127_ _15127_/Q _15127_/CLK _15127_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12339_ VPWR VGND VGND VPWR _12339_/X hold757/A _12339_/B sky130_fd_sc_hd__or2_1
XFILLER_12_1089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_64_1400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15058_ _15058_/Q _15058_/CLK _15058_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_49_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07880_ VGND VPWR VGND VPWR _07668_/B _07813_/A _08104_/B _07880_/X _07311_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_1224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09550_ VGND VPWR VPWR VGND _14512_/D _09550_/A1 _09555_/S hold203/X sky130_fd_sc_hd__mux2_1
X_08501_ VPWR VGND VGND VPWR _09923_/D _08505_/C _09912_/A _08502_/B sky130_fd_sc_hd__o21a_1
X_09481_ VGND VPWR VPWR VGND _14575_/D _09863_/A0 _09482_/S hold461/X sky130_fd_sc_hd__mux2_1
X_08432_ VPWR VGND VGND VPWR _08432_/X _15360_/Q _08486_/B sky130_fd_sc_hd__or2_1
X_08363_ VGND VPWR VPWR VGND _15410_/D hold361/X _08375_/S fanout15/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08294_ _08294_/X _08289_/Y _08292_/X _08293_/X _08294_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07314_ VPWR VGND VPWR VGND _07679_/A _07314_/A _07314_/B sky130_fd_sc_hd__or2_2
X_14008__1125 VPWR VGND VPWR VGND _15380_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_07245_ VPWR VGND VPWR VGND _08116_/A _08117_/A sky130_fd_sc_hd__inv_2
X_07176_ VPWR VGND _07316_/A _07315_/B _15469_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout300 VGND VPWR _10472_/S _10484_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout322 VGND VPWR _11241_/S _11240_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13540__657 VPWR VGND VPWR VGND _14871_/CLK clkload17/A sky130_fd_sc_hd__inv_2
Xfanout311 VGND VPWR _10735_/S _10730_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13937__1054 VPWR VGND VPWR VGND _15309_/CLK clkload31/A sky130_fd_sc_hd__inv_2
Xfanout344 VGND VPWR _10795_/S _11216_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout333 VGND VPWR _11068_/S _11175_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout355 VGND VPWR _08195_/C _10288_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout366 VPWR VGND _10985_/S fanout382/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout388 VPWR VGND _10486_/A1 _10705_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout377 VPWR VGND _10315_/S fanout381/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_47_729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09817_ VGND VPWR VPWR VGND _14235_/D fanout31/X _09833_/S hold185/X sky130_fd_sc_hd__mux2_1
Xfanout399 VGND VPWR _11252_/C1 _11185_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1252 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09748_ VGND VPWR VPWR VGND _14298_/D fanout27/X _09756_/S hold621/X sky130_fd_sc_hd__mux2_1
X_13393__510 VPWR VGND VPWR VGND _14668_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_11710_ VPWR VGND VGND VPWR _11710_/X hold406/A _12716_/S sky130_fd_sc_hd__or2_1
X_09679_ VGND VPWR VPWR VGND _14361_/D hold949/X _09693_/S fanout26/X sky130_fd_sc_hd__mux2_1
X_12690_ VPWR VGND VGND VPWR _12690_/X _12698_/S _12690_/B sky130_fd_sc_hd__or2_1
X_13434__551 VPWR VGND VPWR VGND _14709_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_11641_ VPWR VGND VGND VPWR _11622_/Y _11640_/X _10710_/B _15446_/Q _15446_/D _11296_/A
+ sky130_fd_sc_hd__o221a_1
X_11572_ VPWR VGND VGND VPWR _11572_/X _12098_/A _11572_/B sky130_fd_sc_hd__or2_1
X_14360_ hold857/A _14360_/CLK _14360_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10523_ VGND VPWR VGND VPWR _10523_/X _10520_/X _10522_/X _10523_/A1 _10634_/C1 sky130_fd_sc_hd__a211o_1
X_14291_ hold169/A _14291_/CLK _14291_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10454_ VGND VPWR VPWR VGND _10454_/X _14485_/Q _10464_/S hold545/A sky130_fd_sc_hd__mux2_1
X_10385_ VGND VPWR VPWR VGND _10385_/X _10382_/X _10685_/S _10381_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12124_ VGND VPWR VPWR VGND _12124_/X hold996/A _12149_/S hold533/A sky130_fd_sc_hd__mux2_1
X_12055_ VGND VPWR VPWR VGND _12055_/X _12052_/X _12221_/S _12051_/X sky130_fd_sc_hd__mux2_1
X_11006_ VPWR VGND VPWR VGND _11005_/X _11210_/A _12491_/B1 _11006_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11908_ VPWR VGND VPWR VGND _11907_/X _12212_/A1 _11906_/X _11908_/Y sky130_fd_sc_hd__a21oi_1
X_11839_ VPWR VGND VGND VPWR _11839_/X _12174_/S _11839_/B sky130_fd_sc_hd__or2_1
X_14627_ hold623/A _14627_/CLK _14627_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13177__294 VPWR VGND VPWR VGND _14452_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_14558_ hold490/A _14558_/CLK _14558_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14489_ _14489_/Q _14489_/CLK _14489_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08981_ VGND VPWR VGND VPWR _08981_/X _15478_/Q _08972_/A hold944/X _08980_/Y sky130_fd_sc_hd__a211o_1
X_07932_ VPWR VGND VGND VPWR _07886_/A _07915_/Y _07993_/A _07931_/X _07932_/X sky130_fd_sc_hd__o22a_1
X_12910__27 VPWR VGND VPWR VGND _14152_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_13875__992 VPWR VGND VPWR VGND _15247_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_07863_ VPWR VGND VPWR VGND _07906_/A _15564_/Q _15565_/Q _07864_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_1308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09602_ VGND VPWR VPWR VGND _14466_/D fanout58/X _09619_/S hold716/X sky130_fd_sc_hd__mux2_1
X_07794_ _07992_/B _07727_/X _07794_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_09533_ VGND VPWR VPWR VGND _14529_/D fanout54/X _09549_/S hold168/X sky130_fd_sc_hd__mux2_1
XFILLER_37_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13418__535 VPWR VGND VPWR VGND _14693_/CLK clkload39/A sky130_fd_sc_hd__inv_2
X_09464_ VGND VPWR VPWR VGND _14592_/D clone100/X _09482_/S hold254/X sky130_fd_sc_hd__mux2_1
XFILLER_64_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08415_ VPWR VGND VGND VPWR hold280/A _08415_/B _08415_/Y sky130_fd_sc_hd__nand2b_1
X_09395_ VGND VPWR VPWR VGND _14654_/D _09408_/S hold1119/X clone44/X sky130_fd_sc_hd__mux2_4
XFILLER_19_1029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_75_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08346_ VGND VPWR VPWR VGND _15427_/D hold448/X _08356_/S clone45/A sky130_fd_sc_hd__mux2_1
X_08277_ VGND VPWR VPWR VGND _08277_/X _08276_/Y _08277_/S _08275_/X sky130_fd_sc_hd__mux2_1
X_07228_ VGND VPWR VGND VPWR _08278_/A _07143_/X _07223_/X _14380_/Q _15446_/Q sky130_fd_sc_hd__a211o_1
XFILLER_4_806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07159_ VPWR VGND VPWR VGND _07625_/A _07159_/A _07626_/A sky130_fd_sc_hd__or2_2
X_10170_ VGND VPWR VGND VPWR _10170_/X _14253_/Q _10688_/A2 _10169_/X _10467_/S sky130_fd_sc_hd__o211a_1
X_12985__102 VPWR VGND VPWR VGND _14228_/CLK clkload17/A sky130_fd_sc_hd__inv_2
Xfanout130 VGND VPWR _09548_/A1 _09686_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout152 VPWR VGND VPWR VGND _08540_/A2 _08502_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout141 VPWR VGND _08627_/C1 _08730_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout163 VPWR VGND _08691_/B1 _08522_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout174 VGND VPWR _08298_/A1 _12147_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout185 VGND VPWR _12373_/A _12735_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout196 VGND VPWR _11638_/A1 _12099_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_28_751 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12811_ VGND VPWR VPWR VGND _15560_/D _12810_/Y _12809_/X _12834_/C1 _07544_/X _09975_/A
+ sky130_fd_sc_hd__a32o_1
Xtt_um_femto_890 uio_oe[1] tt_um_femto_890/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_12742_ VPWR VGND VGND VPWR _12742_/X _14998_/Q _12747_/S sky130_fd_sc_hd__or2_1
X_15530_ hold266/A _15530_/CLK _15530_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_69_Right_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15461_ VGND VPWR VGND VPWR _15461_/Q _15461_/D clkload20/A sky130_fd_sc_hd__dfxtp_4
X_12673_ VGND VPWR VGND VPWR _12673_/X _15028_/Q _12743_/A2 _12735_/S _12672_/X sky130_fd_sc_hd__o211a_1
XFILLER_42_286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_31_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11624_ VGND VPWR VPWR VGND _11624_/X hold871/A _12089_/S hold648/A sky130_fd_sc_hd__mux2_1
X_14412_ hold983/A _14412_/CLK _14412_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15392_ hold698/A _15392_/CLK _15392_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11555_ VPWR VGND VGND VPWR _11555_/A _11555_/Y _11555_/B sky130_fd_sc_hd__nand2_1
X_14343_ hold564/A _14343_/CLK _14343_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_633 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11486_ VGND VPWR VPWR VGND _15079_/D _11485_/X _11492_/S hold1417/X sky130_fd_sc_hd__mux2_1
X_12976__93 VPWR VGND VPWR VGND _14219_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_10506_ VGND VPWR VPWR VGND _10507_/B _10505_/Y _10617_/S _10497_/Y sky130_fd_sc_hd__mux2_1
X_13211__328 VPWR VGND VPWR VGND _14486_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_14274_ hold552/A _14274_/CLK _14274_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10437_ VGND VPWR VPWR VGND _10437_/X _14871_/Q _10553_/S hold612/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_78_Right_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_1214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_48_1247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10368_ VGND VPWR VPWR VGND _10368_/X hold486/A _10632_/B hold447/A sky130_fd_sc_hd__mux2_1
X_13859__976 VPWR VGND VPWR VGND _15231_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_2_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10299_ VGND VPWR VGND VPWR _10299_/X hold958/A _10633_/A2 _10298_/X _10510_/S sky130_fd_sc_hd__o211a_1
X_12107_ VPWR VGND VGND VPWR _12107_/X hold430/A _12112_/S sky130_fd_sc_hd__or2_1
XFILLER_61_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12038_ VGND VPWR VPWR VGND _12038_/X hold902/A _12043_/B hold352/A sky130_fd_sc_hd__mux2_1
X_13105__222 VPWR VGND VPWR VGND _14348_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_14007__1124 VPWR VGND VPWR VGND _15379_/CLK clkload16/A sky130_fd_sc_hd__inv_2
XFILLER_22_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08200_ VPWR VGND VGND VPWR _08240_/A _08200_/Y _08200_/B sky130_fd_sc_hd__nand2_1
X_13936__1053 VPWR VGND VPWR VGND _15308_/CLK clkload31/A sky130_fd_sc_hd__inv_2
X_09180_ VGND VPWR VPWR VGND _14911_/D hold466/X _09188_/S fanout36/X sky130_fd_sc_hd__mux2_1
XFILLER_21_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08131_ VGND VPWR VGND VPWR _08252_/A2 _15145_/Q _08132_/A _08130_/X sky130_fd_sc_hd__a21oi_2
X_08062_ VGND VPWR _08066_/A _12790_/B _08062_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13803__920 VPWR VGND VPWR VGND _15175_/CLK clkload13/A sky130_fd_sc_hd__inv_2
XFILLER_31_1284 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08964_ VGND VPWR VGND VPWR _15116_/D hold588/X _08985_/A2 _08963_/X _08955_/A sky130_fd_sc_hd__o211a_1
X_07915_ VGND VPWR _07915_/B _07915_/Y _07915_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_08895_ VGND VPWR VGND VPWR _15145_/D _15144_/Q _08902_/B _08894_/X _11382_/S sky130_fd_sc_hd__o211a_1
XFILLER_57_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07846_ VPWR VGND VGND VPWR _08220_/A _07846_/B _07846_/Y sky130_fd_sc_hd__nor2_1
X_07777_ VPWR VGND VGND VPWR _07777_/A _07777_/B _08210_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09516_ VGND VPWR VPWR VGND _14543_/D _09863_/A0 _09517_/S hold804/X sky130_fd_sc_hd__mux2_1
X_13652__769 VPWR VGND VPWR VGND _14992_/CLK clkload38/A sky130_fd_sc_hd__inv_2
X_09447_ VGND VPWR VPWR VGND _14605_/D _09865_/A0 _09449_/S hold882/X sky130_fd_sc_hd__mux2_1
X_09378_ VGND VPWR VPWR VGND _14668_/D hold702/X _09379_/S _09658_/A0 sky130_fd_sc_hd__mux2_1
X_08329_ VGND VPWR VPWR VGND _15490_/D fanout5/X _08338_/S hold750/X sky130_fd_sc_hd__mux2_1
X_11340_ VPWR VGND VGND VPWR _11340_/A _11340_/B _14832_/D sky130_fd_sc_hd__nor2_1
XFILLER_10_1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11271_ VPWR VGND VGND VPWR _11549_/B _15434_/Q _11271_/B sky130_fd_sc_hd__or2_1
X_13546__663 VPWR VGND VPWR VGND _14877_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_10222_ VGND VPWR VGND VPWR _10222_/X hold997/A _11003_/A2 _10221_/X _10985_/S sky130_fd_sc_hd__o211a_1
X_10153_ VGND VPWR VGND VPWR _10153_/X _10150_/X _10152_/X _10347_/A1 _10608_/A1 sky130_fd_sc_hd__a211o_1
X_14961_ hold738/A _14961_/CLK _14961_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10084_ VGND VPWR VPWR VGND _10084_/X hold897/A _10271_/S hold625/A sky130_fd_sc_hd__mux2_1
X_14892_ _14892_/Q _14892_/CLK _14892_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10986_ VPWR VGND VPWR VGND _10985_/X _11237_/A1 _10984_/X _10986_/Y sky130_fd_sc_hd__a21oi_1
X_15513_ hold192/A _15513_/CLK _15513_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12725_ VGND VPWR VPWR VGND _12725_/X _14218_/Q _12726_/S _15226_/Q sky130_fd_sc_hd__mux2_1
X_15444_ _15444_/Q clkload47/A _15444_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12656_ VPWR VGND VPWR VGND _12655_/X _12656_/A1 _12654_/X _12656_/Y sky130_fd_sc_hd__a21oi_1
X_12587_ VGND VPWR VPWR VGND _12587_/X hold458/A _12599_/S hold354/A sky130_fd_sc_hd__mux2_1
X_11607_ VGND VPWR VPWR VGND _11607_/X hold780/A _11838_/S hold318/A sky130_fd_sc_hd__mux2_1
X_15375_ hold765/A _15375_/CLK _15375_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14326_ hold739/A _14326_/CLK _14326_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11538_ VGND VPWR VPWR VGND _15096_/D _11537_/X _11538_/S hold1406/X sky130_fd_sc_hd__mux2_1
Xhold408 hold408/X hold408/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ _14257_/Q _14257_/CLK _14257_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold419 hold419/X hold419/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ VGND VPWR VPWR VGND _11469_/X _15075_/Q _11475_/S _15073_/Q sky130_fd_sc_hd__mux2_1
X_14188_ _14188_/Q _14188_/CLK _14188_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1108 hold1108/X _15346_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 hold1119/X _14654_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ VGND VPWR VGND VPWR _07700_/X _08002_/B1 _07692_/Y _15594_/Q _07699_/X sky130_fd_sc_hd__a211o_1
X_08680_ VGND VPWR VGND VPWR _15288_/D hold890/X _08686_/A2 _08679_/X _12492_/C1 sky130_fd_sc_hd__o211a_1
X_07631_ VGND VPWR VGND VPWR _07631_/X _15133_/Q _15360_/Q clone13/X _08034_/B1 sky130_fd_sc_hd__a22o_4
XFILLER_54_827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07562_ VPWR VGND VPWR VGND _12878_/A _07827_/D _15572_/Q _07563_/B sky130_fd_sc_hd__or3_1
XFILLER_4_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09301_ VGND VPWR VPWR VGND _14740_/D fanout6/X _09302_/S hold312/X sky130_fd_sc_hd__mux2_1
X_13489__606 VPWR VGND VPWR VGND _14764_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_07493_ VGND VPWR VPWR VGND _15453_/Q _08592_/B _15598_/Q sky130_fd_sc_hd__xor2_1
X_09232_ VPWR VGND VPWR VGND _08413_/Y _09239_/B _09938_/A _09232_/B sky130_fd_sc_hd__or3b_2
XFILLER_72_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09163_ VGND VPWR VPWR VGND _14935_/D fanout96/X _09163_/S hold922/X sky130_fd_sc_hd__mux2_1
X_08114_ VPWR VGND VPWR VGND _11440_/B _08113_/X _08114_/Y _07331_/A _08112_/A sky130_fd_sc_hd__a22oi_1
X_13233__350 VPWR VGND VPWR VGND _14508_/CLK clkload6/A sky130_fd_sc_hd__inv_2
XFILLER_68_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09094_ VGND VPWR VPWR VGND _14999_/D hold1086/X _09094_/S fanout96/X sky130_fd_sc_hd__mux2_1
Xhold920 hold920/X hold920/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08045_ VPWR VGND VGND VPWR _08240_/A _10064_/C _08045_/Y sky130_fd_sc_hd__nor2_1
Xhold931 hold931/X hold931/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 hold942/X hold942/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 hold953/X hold953/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold964 hold964/X hold964/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 hold986/X hold986/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 hold975/X hold975/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 hold997/X hold997/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ VGND VPWR _10000_/B _15614_/Q _15613_/Q _09996_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_08947_ VPWR VGND _15124_/D _08947_/B _11567_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_76_429 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08878_ VPWR VGND VGND VPWR _08878_/X _15153_/Q _08926_/B sky130_fd_sc_hd__or2_1
XFILLER_28_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13082__199 VPWR VGND VPWR VGND _14325_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_07829_ VGND VPWR VGND VPWR _12817_/A _10078_/A _12833_/A sky130_fd_sc_hd__or2_4
X_10840_ VGND VPWR VPWR VGND _10840_/X hold880/A _10850_/S hold652/A sky130_fd_sc_hd__mux2_1
XFILLER_60_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_25_540 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10771_ VGND VPWR VGND VPWR _10771_/X hold808/A _11262_/A2 _10770_/X _11215_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_25_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12510_ VPWR VGND VGND VPWR _12658_/A _12510_/B _12510_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12441_ VGND VPWR VGND VPWR _12441_/X hold961/A _12669_/A2 _12662_/A1 _12440_/X sky130_fd_sc_hd__o211a_1
XFILLER_51_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14006__1123 VPWR VGND VPWR VGND _15378_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_15160_ _15160_/Q _15160_/CLK _15160_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12372_ VGND VPWR VPWR VGND _12372_/X _15387_/Q _12372_/S _15534_/Q sky130_fd_sc_hd__mux2_1
X_11323_ VPWR VGND _14826_/D _11323_/B _11327_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_12946__63 VPWR VGND VPWR VGND _14189_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_13780__897 VPWR VGND VPWR VGND _15152_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_15091_ _15091_/Q clkload33/A _15091_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11254_ VGND VPWR VGND VPWR _11254_/X _11253_/X _11252_/X _11250_/S _11254_/C1 sky130_fd_sc_hd__a211o_1
X_10205_ VGND VPWR VPWR VGND _10205_/X hold937/A _10567_/S hold423/A sky130_fd_sc_hd__mux2_1
XFILLER_4_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11185_ VGND VPWR VGND VPWR _11185_/X _11182_/X _11184_/X _11185_/A1 _11185_/C1 sky130_fd_sc_hd__a211o_1
X_13935__1052 VPWR VGND VPWR VGND _15307_/CLK clkload31/A sky130_fd_sc_hd__inv_2
XFILLER_48_621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10136_ VGND VPWR VPWR VGND _10137_/B _10135_/Y _10617_/S _10127_/Y sky130_fd_sc_hd__mux2_1
X_10067_ VPWR VGND VGND VPWR _07665_/Y _07637_/B _07637_/A _07652_/B _10067_/X sky130_fd_sc_hd__o22a_1
X_14944_ hold525/A _14944_/CLK _14944_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14875_ _14875_/Q _14875_/CLK _14875_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13674__791 VPWR VGND VPWR VGND _15014_/CLK clkload11/A sky130_fd_sc_hd__inv_2
XFILLER_21_1250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10969_ VPWR VGND VPWR VGND _10968_/X _11247_/A _12713_/B1 _10969_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_1379 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12708_ VGND VPWR VPWR VGND _12708_/X hold841/A _12708_/S hold509/A sky130_fd_sc_hd__mux2_1
X_13217__334 VPWR VGND VPWR VGND _14492_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_15427_ hold448/A _15427_/CLK _15427_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12639_ VPWR VGND VPWR VGND _12638_/X _12658_/A _12713_/B1 _12639_/X sky130_fd_sc_hd__a21o_1
X_15358_ _15358_/Q _15358_/CLK _15358_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14309_ hold373/A _14309_/CLK _14309_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15289_ _15289_/Q _15289_/CLK _15289_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold205 hold205/X hold205/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 hold216/X hold216/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/X hold249/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/X hold227/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/X hold238/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout707 VGND VPWR _08424_/Y _08488_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout729 VPWR VGND _10192_/B _10562_/B VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_63_1339 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout718 VGND VPWR _10056_/Y _12807_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09850_ VGND VPWR VPWR VGND _14172_/D hold422/X _09865_/S fanout36/X sky130_fd_sc_hd__mux2_1
X_08801_ VGND VPWR VPWR VGND _15208_/D fanout20/X _08806_/S hold181/X sky130_fd_sc_hd__mux2_1
X_09781_ VGND VPWR VPWR VGND _14268_/D fanout35/X _09790_/S hold544/X sky130_fd_sc_hd__mux2_1
X_08732_ VPWR VGND VPWR VGND _15264_/Q _15266_/Q _15267_/Q _15265_/Q _08853_/A sky130_fd_sc_hd__or4_1
X_08663_ VGND VPWR VGND VPWR _15293_/D hold883/X _08704_/A2 _08662_/X _08717_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_22_1058 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08594_ VPWR VGND VGND VPWR _08617_/A _08995_/B _08594_/Y sky130_fd_sc_hd__nor2_1
X_07614_ VPWR VGND VPWR VGND _07614_/B _07614_/C _07614_/A _07614_/X sky130_fd_sc_hd__or3_4
X_07545_ VGND VPWR _07545_/B _07545_/Y _07545_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07476_ VPWR VGND VGND VPWR _15446_/Q _07476_/Y _07476_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09215_ VGND VPWR VPWR VGND _14878_/D hold1026/X _09229_/S fanout31/X sky130_fd_sc_hd__mux2_1
X_09146_ VGND VPWR VPWR VGND _14952_/D fanout35/X _09161_/S hold792/X sky130_fd_sc_hd__mux2_1
XFILLER_30_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09077_ VGND VPWR VPWR VGND _15016_/D hold1082/X _09092_/S fanout37/X sky130_fd_sc_hd__mux2_1
X_08028_ VPWR VGND VGND VPWR _08028_/A _08104_/B _08028_/Y sky130_fd_sc_hd__nor2_1
X_13010__127 VPWR VGND VPWR VGND _14253_/CLK clkload24/A sky130_fd_sc_hd__inv_2
Xhold761 hold761/X hold761/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_1_414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold772 hold772/X hold772/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 hold750/X hold750/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 hold794/X hold794/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 hold783/X hold783/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09979_ VGND VPWR VGND VPWR _09979_/X _08425_/A _15365_/Q _14767_/Q sky130_fd_sc_hd__a21bo_1
XFILLER_79_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1461 _07102_/A _15347_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13658__775 VPWR VGND VPWR VGND _14998_/CLK clkload49/A sky130_fd_sc_hd__inv_2
Xhold1450 hold1450/X _15295_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11941_ VGND VPWR VGND VPWR _11941_/X _11938_/X _11940_/X _11968_/S _12175_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_18_838 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11872_ VGND VPWR VPWR VGND _11872_/X _14195_/Q _11876_/B hold252/A sky130_fd_sc_hd__mux2_1
X_14660_ hold592/A _14660_/CLK _14660_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10823_ VGND VPWR VPWR VGND _10823_/X hold720/A _11091_/S hold741/A sky130_fd_sc_hd__mux2_1
X_14591_ hold526/A _14591_/CLK _14591_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_44_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_1043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10754_ VGND VPWR VGND VPWR _10754_/X _11086_/C1 _10750_/X _10753_/X _11217_/C1 sky130_fd_sc_hd__o211a_1
X_10685_ VGND VPWR VPWR VGND _10685_/X _10684_/X _10685_/S _10683_/X sky130_fd_sc_hd__mux2_1
X_12424_ VGND VPWR VGND VPWR _12424_/X _12662_/A1 _12420_/X _12423_/X _12662_/C1 sky130_fd_sc_hd__o211a_1
X_15212_ hold550/A _15212_/CLK _15212_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12355_ VGND VPWR VPWR VGND _12355_/X _12354_/X _12367_/S _12353_/X sky130_fd_sc_hd__mux2_1
X_15143_ _15143_/Q _15143_/CLK _15143_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11306_ VGND VPWR VGND VPWR _14820_/D _14381_/Q _11303_/B _11305_/X _11308_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_5_764 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12286_ VPWR VGND VPWR VGND _12285_/X _12703_/A1 _12284_/X _12286_/Y sky130_fd_sc_hd__a21oi_1
X_15074_ _15074_/Q clkload14/A _15074_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11237_ VPWR VGND VPWR VGND _11236_/X _11237_/A1 _11235_/X _11237_/Y sky130_fd_sc_hd__a21oi_1
X_11168_ VPWR VGND VGND VPWR _11168_/X _11170_/S _11168_/B sky130_fd_sc_hd__or2_1
X_10119_ VPWR VGND VGND VPWR _10100_/Y _10118_/X _10710_/B _14379_/Q _14379_/D _11296_/A
+ sky130_fd_sc_hd__o221a_1
X_11099_ VGND VPWR VPWR VGND _11099_/X _14374_/Q _11109_/S _14726_/Q sky130_fd_sc_hd__mux2_1
XFILLER_48_440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_23_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14927_ _14927_/Q clkload28/A _14927_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14858_ _14858_/Q clkload26/A _14858_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14789_ _14789_/Q _14789_/CLK _14789_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07330_ VPWR VGND VGND VPWR _07574_/A _08286_/B _07331_/A sky130_fd_sc_hd__nor2_4
X_13451__568 VPWR VGND VPWR VGND _14726_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_09000_ VGND VPWR VGND VPWR _09000_/X hold1125/X _09015_/A2 _08999_/X _09000_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07261_ VPWR VGND VGND VPWR _14394_/Q _07230_/S _07265_/B1 _07263_/B sky130_fd_sc_hd__o21a_1
Xclkbuf_3_7_0_clk clkload5/A clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07192_ VPWR VGND _07195_/A _07355_/B _15455_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_09902_ VPWR VGND VPWR VGND _09900_/A _15480_/Q _09907_/S _09902_/X sky130_fd_sc_hd__a21o_1
Xfanout515 VGND VPWR _12372_/S _12370_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13345__462 VPWR VGND VPWR VGND _14620_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
Xfanout504 VPWR VGND _12220_/S _12227_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout537 VGND VPWR fanout538/X _12577_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout548 VPWR VGND _08495_/A2 clone13/A VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout526 VGND VPWR fanout539/X _12446_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09833_ VGND VPWR VPWR VGND _14219_/D fanout97/X _09833_/S hold320/X sky130_fd_sc_hd__mux2_1
Xfanout559 VPWR VGND _09721_/S _09694_/Y VPWR VGND sky130_fd_sc_hd__buf_4
X_09764_ VPWR VGND VGND VPWR _09799_/B _09764_/Y _09764_/A sky130_fd_sc_hd__nor2_2
XFILLER_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_473 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08715_ VGND VPWR VGND VPWR _15276_/D hold982/X _08721_/A2 _08714_/X _08717_/C1 sky130_fd_sc_hd__o211a_1
X_09695_ VPWR VGND VPWR VGND _09695_/Y _09725_/S sky130_fd_sc_hd__inv_2
X_14005__1122 VPWR VGND VPWR VGND _15377_/CLK clkload11/A sky130_fd_sc_hd__inv_2
Xrebuffer42 VPWR VGND VPWR VGND rebuffer42/X rebuffer43/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_55_966 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer31 VPWR VGND VPWR VGND rebuffer31/X rebuffer32/X sky130_fd_sc_hd__dlygate4sd1_1
X_08646_ VPWR VGND VGND VPWR _08645_/X _08690_/S _08194_/Y _14407_/Q _08646_/X _08644_/X
+ sky130_fd_sc_hd__o221a_1
X_08577_ VPWR VGND VGND VPWR _08582_/A _08986_/B _08577_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_1287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07528_ VPWR VGND VPWR VGND _07551_/A _07551_/B _07530_/A _07506_/A _07433_/A sky130_fd_sc_hd__a211oi_2
X_07459_ VPWR VGND VGND VPWR _08597_/B _15452_/Q _15597_/Q sky130_fd_sc_hd__or2_1
XFILLER_50_693 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13934__1051 VPWR VGND VPWR VGND _15306_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_10470_ VPWR VGND VGND VPWR _10507_/A _10470_/B _10470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_517 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09129_ VPWR VGND VGND VPWR _09694_/A _09129_/Y _09198_/C sky130_fd_sc_hd__nor2_2
X_12916__33 VPWR VGND VPWR VGND _14159_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_12140_ VPWR VGND VGND VPWR _12214_/A _12140_/B _12140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold580 hold580/X hold580/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12071_ VGND VPWR VGND VPWR _12071_/X hold894/A _12080_/A2 _12230_/A1 _12070_/X sky130_fd_sc_hd__o211a_1
XFILLER_46_1367 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11022_ VGND VPWR VPWR VGND _11022_/X _11019_/X _11162_/S _11018_/X sky130_fd_sc_hd__mux2_1
Xhold591 hold591/X hold591/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1280 _08734_/B _15262_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1291 _15344_/D _08465_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14209__927 _14209_/D _14209__927/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_14712_ hold634/A _14712_/CLK _14712_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_17_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11924_ VGND VPWR VPWR VGND _11924_/X hold981/A _12149_/S hold674/A sky130_fd_sc_hd__mux2_1
X_14643_ hold443/A _14643_/CLK _14643_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11855_ VGND VPWR VGND VPWR _11855_/X _15006_/Q _12040_/A2 _12174_/S _11854_/X sky130_fd_sc_hd__o211a_1
X_10806_ VGND VPWR VPWR VGND _10806_/X hold743/A _11216_/S hold585/A sky130_fd_sc_hd__mux2_1
X_14574_ hold219/A _14574_/CLK _14574_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11786_ VGND VPWR VGND VPWR _11786_/X _11783_/X _11785_/X _12008_/A1 _12008_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_9_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10737_ VGND VPWR VGND VPWR _10737_/X _10745_/C1 _10732_/X _10736_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_13288__405 VPWR VGND VPWR VGND _14563_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_10668_ VPWR VGND VGND VPWR _10668_/X hold241/A _10670_/S sky130_fd_sc_hd__or2_1
X_12407_ VGND VPWR VGND VPWR _12407_/X _12415_/C1 _12402_/X _12406_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_16_1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10599_ VPWR VGND VPWR VGND _10598_/X _10729_/A _11973_/B _10599_/X sky130_fd_sc_hd__a21o_1
X_15126_ _15126_/Q _15126_/CLK _15126_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12338_ VGND VPWR VPWR VGND _12338_/X hold501/A _12594_/B hold518/A sky130_fd_sc_hd__mux2_1
X_13329__446 VPWR VGND VPWR VGND _14604_/CLK clkload8/A sky130_fd_sc_hd__inv_2
XFILLER_64_1412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12269_ VPWR VGND VGND VPWR _12269_/X _15463_/Q _12269_/B sky130_fd_sc_hd__or2_1
X_15057_ hold385/A _15057_/CLK _15057_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08500_ VPWR VGND VPWR VGND _08500_/B _08500_/C hold239/A _08505_/C _14140_/Q sky130_fd_sc_hd__or4b_1
X_09480_ VGND VPWR VPWR VGND _14576_/D _09723_/A1 _09485_/S hold195/X sky130_fd_sc_hd__mux2_1
XFILLER_64_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08431_ VGND VPWR VGND VPWR _15361_/D hold1367/X _08485_/A2 _08430_/X _11388_/S sky130_fd_sc_hd__o211a_1
XFILLER_37_999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_37_988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08362_ VGND VPWR VPWR VGND _15411_/D hold437/X _08366_/S fanout19/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08293_ VGND VPWR VPWR VGND _08293_/X _08293_/A3 _08290_/B _15445_/Q _08293_/B1 _15065_/Q
+ sky130_fd_sc_hd__a32o_1
X_07313_ VPWR VGND VGND VPWR _07313_/A _07693_/A _07313_/B sky130_fd_sc_hd__nand2_1
X_07244_ VPWR VGND VGND VPWR _07244_/A _08117_/A _07244_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_1345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07175_ VPWR VGND VGND VPWR _14403_/Q _07301_/A2 _07301_/B1 _07315_/B sky130_fd_sc_hd__o21a_1
Xfanout301 VPWR VGND _10472_/S fanout314/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout323 VGND VPWR _11102_/S _11109_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout312 VGND VPWR _10742_/S _10735_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout345 VGND VPWR _11093_/S _11091_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_59_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout356 VGND VPWR _10677_/S _10685_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout334 VGND VPWR _11068_/S _11165_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_59_568 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout389 VPWR VGND _10705_/A fanout390/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout378 VGND VPWR _11205_/A _11213_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_47_708 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09816_ VGND VPWR VPWR VGND _14236_/D fanout35/X _09825_/S hold334/X sky130_fd_sc_hd__mux2_1
Xfanout367 VGND VPWR _11244_/S _10911_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13122__239 VPWR VGND VPWR VGND _14365_/CLK _12962__79/A sky130_fd_sc_hd__inv_2
X_09747_ VGND VPWR VPWR VGND _14299_/D fanout31/X _09763_/S hold196/X sky130_fd_sc_hd__mux2_1
XFILLER_36_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_55_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_936 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09678_ VGND VPWR VPWR VGND _14362_/D hold918/X _09684_/S _08014_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_947 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08629_ VGND VPWR VGND VPWR _08700_/A2 _14386_/Q _08194_/B _08629_/X sky130_fd_sc_hd__o21ba_1
X_11640_ VPWR VGND VPWR VGND _11639_/X _12103_/A _12121_/B1 _11640_/X sky130_fd_sc_hd__a21o_1
X_13473__590 VPWR VGND VPWR VGND _14748_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_11571_ VGND VPWR VPWR VGND _11571_/X hold803/A _11756_/S hold199/A sky130_fd_sc_hd__mux2_1
X_10522_ VGND VPWR VGND VPWR _10522_/X _15010_/Q _10633_/A2 _10521_/X _10510_/S sky130_fd_sc_hd__o211a_1
X_13016__133 VPWR VGND VPWR VGND _14259_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_14290_ hold431/A _14290_/CLK _14290_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10453_ VGND VPWR VPWR VGND _10457_/B hold554/A _10464_/S hold607/A sky130_fd_sc_hd__mux2_1
X_10384_ VGND VPWR VGND VPWR _10384_/X _10698_/A1 _10380_/X _10383_/X _10697_/B1 sky130_fd_sc_hd__o211a_1
X_13820__937 VPWR VGND VPWR VGND _15192_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XFILLER_48_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12123_ VGND VPWR VPWR VGND _12127_/B hold515/A _12155_/S hold676/A sky130_fd_sc_hd__mux2_1
XFILLER_78_800 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12054_ VGND VPWR VGND VPWR _12054_/X _12230_/A1 _12050_/X _12053_/X _12226_/C1 sky130_fd_sc_hd__o211a_1
X_11005_ VPWR VGND _11005_/X _11004_/X _11000_/X _10987_/S _10996_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_13714__831 VPWR VGND VPWR VGND _15054_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_11907_ VGND VPWR VPWR VGND _11907_/X _11904_/X _12147_/S _11903_/X sky130_fd_sc_hd__mux2_1
X_11838_ VGND VPWR VPWR VGND _11838_/X _14450_/Q _11838_/S hold282/A sky130_fd_sc_hd__mux2_1
X_14626_ hold567/A _14626_/CLK _14626_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14557_ hold479/A _14557_/CLK _14557_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_40_clk clkload55/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_11769_ VGND VPWR VPWR VGND _11770_/B _11768_/Y _12102_/S _11760_/Y sky130_fd_sc_hd__mux2_1
X_14488_ hold906/A _14488_/CLK _14488_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14004__1121 VPWR VGND VPWR VGND _15376_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_6_881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15109_ hold944/A _15109_/CLK hold945/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08980_ VPWR VGND VGND VPWR _08983_/A _08980_/B _08980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07931_ VPWR VGND VGND VPWR _07931_/X _07931_/A _07931_/B sky130_fd_sc_hd__or2_1
X_07862_ _07870_/B _07858_/X _07859_/Y _07861_/X _08249_/B2 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_13933__1050 VPWR VGND VPWR VGND _15305_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_09601_ VGND VPWR VPWR VGND _14467_/D fanout60/X _09622_/S hold597/X sky130_fd_sc_hd__mux2_1
X_07793_ VPWR VGND _07958_/B _07730_/B _07794_/B _15558_/Q _07727_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_37_741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09532_ VGND VPWR VPWR VGND _14530_/D fanout56/X _09549_/S hold156/X sky130_fd_sc_hd__mux2_1
X_13457__574 VPWR VGND VPWR VGND _14732_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_09463_ VGND VPWR VPWR VGND _14593_/D _09482_/S fanout52/X hold1151/X sky130_fd_sc_hd__mux2_4
X_08414_ hold154/A _14810_/Q hold153/X _09232_/B _08735_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09394_ VGND VPWR VPWR VGND _14655_/D hold741/X _09408_/S fanout46/X sky130_fd_sc_hd__mux2_1
XFILLER_40_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_1393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08345_ VGND VPWR VPWR VGND _15428_/D hold463/X _08356_/S fanout83/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_clk clkload47/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_22_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08276_ VGND VPWR _08276_/B _08276_/Y _10061_/B VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07227_ VGND VPWR VGND VPWR _07229_/A _07143_/X _07224_/X _07110_/Y _07360_/A sky130_fd_sc_hd__a211o_1
X_07158_ VPWR VGND VPWR VGND _07158_/Y _07626_/A sky130_fd_sc_hd__inv_2
X_07089_ VPWR VGND VPWR VGND _11973_/A _15455_/Q sky130_fd_sc_hd__inv_2
Xfanout131 VGND VPWR _08170_/X _09548_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout120 VGND VPWR _08230_/X _09655_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout142 VPWR VGND _08730_/B1 _08508_/X VPWR VGND sky130_fd_sc_hd__buf_4
Xfanout153 VPWR VGND _09016_/B1 _08937_/Y VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_47_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout164 VPWR VGND _12098_/A _11625_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout175 VGND VPWR _08298_/A1 _11925_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout197 VGND VPWR _11638_/A1 _12008_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout186 VGND VPWR _12536_/S _12655_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_12810_ VPWR VGND VGND VPWR _12817_/A _12810_/Y _12810_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_41_1094 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xtt_um_femto_891 uio_oe[2] tt_um_femto_891/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_12741_ VGND VPWR VPWR VGND _12741_/X _15194_/Q _12747_/S _15062_/Q sky130_fd_sc_hd__mux2_1
X_15460_ VGND VPWR VGND VPWR _15460_/Q _15460_/D clkload18/A sky130_fd_sc_hd__dfxtp_4
X_12672_ VPWR VGND VGND VPWR _12672_/X hold340/A _12736_/B sky130_fd_sc_hd__or2_1
X_14411_ hold878/A _14411_/CLK _14411_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11623_ VGND VPWR VPWR VGND _11623_/X hold983/A _12089_/S hold702/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_clk clkload29/A clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_15391_ hold627/A _15391_/CLK _15391_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_23_490 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11554_ VPWR VGND VPWR VGND hold1160/X _11555_/B _11341_/Y _15437_/D sky130_fd_sc_hd__a21oi_1
X_14342_ _14342_/Q _14342_/CLK _14342_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13250__367 VPWR VGND VPWR VGND _14525_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_11485_ VGND VPWR VPWR VGND _11485_/X _11484_/X _11491_/S _15459_/Q sky130_fd_sc_hd__mux2_1
X_14273_ _14273_/Q _14273_/CLK _14273_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10505_ VPWR VGND VPWR VGND _10504_/X _10505_/A1 _10503_/X _10505_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10436_ VGND VPWR VPWR VGND _10436_/X hold525/A _10553_/S hold644/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10367_ VGND VPWR VGND VPWR _10367_/X _10616_/A1 _10362_/X _10366_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_3_862 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10298_ VPWR VGND VGND VPWR _10298_/X hold203/A _10521_/B sky130_fd_sc_hd__or2_1
X_12106_ VGND VPWR VPWR VGND _12106_/X _12105_/X _12106_/S _12104_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12037_ VGND VPWR VGND VPWR _12037_/X _12193_/C1 _12032_/X _12036_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
X_13144__261 VPWR VGND VPWR VGND _14419_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_34_744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14609_ hold374/A _14609_/CLK _14609_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08130_ VPWR VGND VPWR VGND _11302_/A _15340_/Q _08253_/A2 _08130_/X _14824_/Q sky130_fd_sc_hd__a22o_1
X_15589_ _15589_/Q clkload49/A _15589_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_clk _12954__71/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_08061_ VPWR VGND VPWR VGND _15618_/Q _08299_/A2 _08070_/C _07426_/X _08286_/B _08060_/Y
+ sky130_fd_sc_hd__a221o_1
X_08963_ VPWR VGND VGND VPWR _08963_/X _08969_/A _08963_/B sky130_fd_sc_hd__or2_1
X_07914_ VGND VPWR VGND VPWR _07913_/Y _08286_/A _07933_/C _07914_/B1 sky130_fd_sc_hd__a21oi_2
X_08894_ VPWR VGND VGND VPWR _08894_/X _15145_/Q _08924_/B sky130_fd_sc_hd__or2_1
XFILLER_57_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07845_ VGND VPWR _07864_/A _07846_/B _15566_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07776_ VPWR VGND VPWR VGND _07757_/C _15595_/Q _15548_/Q _07777_/B sky130_fd_sc_hd__a21oi_1
Xclone5 VGND VPWR clone5/A clone5/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_37_593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09515_ VGND VPWR VPWR VGND _14544_/D _09723_/A1 _09520_/S hold586/X sky130_fd_sc_hd__mux2_1
X_09446_ VGND VPWR VPWR VGND _14606_/D _09864_/A0 _09446_/S hold368/X sky130_fd_sc_hd__mux2_1
XFILLER_40_725 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09377_ VGND VPWR VPWR VGND _14669_/D hold477/X _09377_/S _09691_/A0 sky130_fd_sc_hd__mux2_1
X_08328_ VGND VPWR VPWR VGND _15491_/D fanout10/X _08330_/S hold1134/X sky130_fd_sc_hd__mux2_1
X_08259_ VGND VPWR _08258_/X _08182_/S _08259_/Y _07362_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
X_11270_ VPWR VGND VGND VPWR _11271_/B _15433_/Q _11545_/B sky130_fd_sc_hd__or2_1
X_13087__204 VPWR VGND VPWR VGND _14330_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_10221_ VPWR VGND VGND VPWR _10221_/X hold275/A _11231_/S sky130_fd_sc_hd__or2_1
X_10152_ VGND VPWR VGND VPWR _10152_/X _15000_/Q _10629_/A2 _10151_/X _10615_/S sky130_fd_sc_hd__o211a_1
X_14960_ hold845/A _14960_/CLK _14960_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10083_ VGND VPWR VPWR VGND _10087_/B hold876/A _10271_/S hold692/A sky130_fd_sc_hd__mux2_1
X_13128__245 VPWR VGND VPWR VGND _14371_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
XFILLER_48_869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14891_ _14891_/Q _14891_/CLK _14891_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14003__1120 VPWR VGND VPWR VGND _15375_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_15512_ _15512_/Q _15512_/CLK _15512_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12724_ VGND VPWR VPWR VGND _12724_/X _14282_/Q _12736_/B _14314_/Q sky130_fd_sc_hd__mux2_1
X_10985_ VGND VPWR VPWR VGND _10985_/X _10982_/X _10985_/S _10981_/X sky130_fd_sc_hd__mux2_1
X_13785__902 VPWR VGND VPWR VGND _15157_/CLK clkload28/A sky130_fd_sc_hd__inv_2
XFILLER_15_276 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15443_ _15443_/Q clkload47/A _15443_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12655_ VGND VPWR VPWR VGND _12655_/X _12652_/X _12655_/S _12651_/X sky130_fd_sc_hd__mux2_1
X_12586_ VGND VPWR VGND VPWR _12586_/X _14889_/Q _12746_/A2 _12591_/S _12585_/X sky130_fd_sc_hd__o211a_1
X_15374_ hold680/A _15374_/CLK _15374_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11606_ VGND VPWR VPWR VGND _11606_/X _14476_/Q _12097_/S hold396/A sky130_fd_sc_hd__mux2_1
X_14325_ hold717/A _14325_/CLK _14325_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11537_ VGND VPWR VPWR VGND _11537_/X _11536_/X _11537_/S _15476_/Q sky130_fd_sc_hd__mux2_1
X_13826__943 VPWR VGND VPWR VGND _15198_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
XFILLER_8_965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold409 hold409/X hold409/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11468_ VGND VPWR VPWR VGND _15073_/D _11467_/X _11477_/S _15073_/Q sky130_fd_sc_hd__mux2_1
X_14256_ hold394/A _14256_/CLK _14256_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11399_ VPWR VGND VPWR VGND _11362_/X _11399_/A1 _11367_/D _11400_/B sky130_fd_sc_hd__a21o_1
X_14187_ _14187_/Q _14187_/CLK _14187_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10419_ VPWR VGND VGND VPWR _10419_/X hold496/A _10720_/S sky130_fd_sc_hd__or2_1
Xhold1109 hold1109/X _15534_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clkload7/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07630_ VGND VPWR VPWR VGND _15542_/D fanout80/X _08231_/S hold294/X sky130_fd_sc_hd__mux2_1
X_07561_ VPWR VGND VPWR VGND _15136_/Q _08252_/A2 _15363_/Q _08253_/A2 _07561_/X sky130_fd_sc_hd__a22o_2
XFILLER_4_1194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09300_ VGND VPWR VPWR VGND _14741_/D fanout8/X _09310_/S hold304/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07492_ VPWR VGND VGND VPWR _07492_/A _07492_/B _08592_/A sky130_fd_sc_hd__nor2_1
X_09231_ VGND VPWR VPWR VGND _14862_/D hold860/X _09231_/S fanout95/X sky130_fd_sc_hd__mux2_1
XFILLER_72_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09162_ VGND VPWR VPWR VGND _14936_/D _09692_/A0 _09163_/S hold873/X sky130_fd_sc_hd__mux2_1
X_13569__686 VPWR VGND VPWR VGND _14900_/CLK clkload55/A sky130_fd_sc_hd__inv_2
X_08113_ VGND VPWR VPWR VGND _08113_/X _08112_/A _08195_/A _07676_/A sky130_fd_sc_hd__mux2_1
X_09093_ VGND VPWR VPWR VGND _15000_/D hold1112/X _09094_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
Xhold921 hold921/X hold921/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold910 hold910/X hold910/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08044_ VGND VPWR _08044_/B _10064_/C _08047_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold954 hold954/X hold954/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 hold932/X hold932/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 hold943/X hold943/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 hold976/X hold976/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 hold998/X hold998/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 hold965/X hold965/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold987 hold987/X hold987/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09995_ VGND VPWR VPWR VGND _09995_/A _15613_/D _09996_/C sky130_fd_sc_hd__xor2_1
X_08946_ VPWR VGND VPWR VGND _08972_/A _15123_/Q _08933_/A _08947_/B hold1423/X sky130_fd_sc_hd__a22o_1
XFILLER_44_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_28_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08877_ VGND VPWR VGND VPWR _08877_/X hold1249/X _08919_/A2 _08876_/X _11308_/C1
+ sky130_fd_sc_hd__o211a_1
X_07828_ VPWR VGND VGND VPWR _10078_/A _12817_/A _07828_/Y sky130_fd_sc_hd__nor2_1
X_07759_ VPWR VGND _07759_/X _07760_/B _15547_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_44_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10770_ VPWR VGND VGND VPWR _10770_/X hold581/A _11091_/S sky130_fd_sc_hd__or2_1
XFILLER_40_500 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09429_ VGND VPWR VPWR VGND _14623_/D fanout46/X _09443_/S hold720/X sky130_fd_sc_hd__mux2_1
X_13513__630 VPWR VGND VPWR VGND _14788_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_12440_ VPWR VGND VGND VPWR _12440_/X hold834/A _12623_/S sky130_fd_sc_hd__or2_1
XFILLER_40_599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_12_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12371_ VGND VPWR VPWR VGND _12371_/X _15502_/Q _12599_/S _14528_/Q sky130_fd_sc_hd__mux2_1
X_11322_ VGND VPWR VPWR VGND _11323_/B _11342_/C _11320_/Y _11313_/C _11317_/X _14826_/Q
+ sky130_fd_sc_hd__a32o_1
X_15090_ _15090_/Q clkload33/A _15090_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13912__1029 VPWR VGND VPWR VGND _15284_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_11253_ VGND VPWR VPWR VGND _11253_/X _14893_/Q _11261_/B _15429_/Q sky130_fd_sc_hd__mux2_1
XFILLER_45_1207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10204_ VGND VPWR VPWR VGND _10204_/X _14190_/Q _10994_/S hold190/A sky130_fd_sc_hd__mux2_1
X_12961__78 VPWR VGND VPWR VGND _14204_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_11184_ VGND VPWR VGND VPWR _11184_/X hold959/A _11184_/A2 _11183_/X _11250_/S sky130_fd_sc_hd__o211a_1
X_13362__479 VPWR VGND VPWR VGND _14637_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_10135_ VPWR VGND VPWR VGND _10134_/X _10616_/A1 _10133_/X _10135_/Y sky130_fd_sc_hd__a21oi_1
X_14943_ hold835/A _14943_/CLK _14943_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10066_ VPWR VGND VGND VPWR _10065_/X _10066_/C _10066_/Y _10066_/B _10066_/A sky130_fd_sc_hd__nor4b_1
X_14874_ _14874_/Q _14874_/CLK _14874_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10968_ VPWR VGND _10968_/X _10967_/X _10963_/X _11246_/S _10959_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_43_393 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12707_ VGND VPWR VGND VPWR _12707_/X _12706_/X _12705_/X _11810_/S _12748_/C1 sky130_fd_sc_hd__a211o_1
X_13256__373 VPWR VGND VPWR VGND _14531_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_28_Left_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10899_ VGND VPWR VPWR VGND _10899_/X _14337_/Q _10919_/S _15249_/Q sky130_fd_sc_hd__mux2_1
X_15426_ hold363/A _15426_/CLK _15426_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12638_ VPWR VGND _12638_/X _12637_/X _12633_/X _12731_/S _12629_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12569_ VGND VPWR VPWR VGND _12569_/X _14342_/Q _12577_/S _15254_/Q sky130_fd_sc_hd__mux2_1
X_15357_ _15357_/Q _15357_/CLK _15357_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold217 hold217/X hold217/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 hold206/X hold206/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ hold890/A _15288_/CLK _15288_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14308_ hold370/A _14308_/CLK _14308_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold239 hold239/X hold239/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_1421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14239_ hold244/A _14239_/CLK _14239_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold228 hold228/X hold228/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout708 VGND VPWR _08486_/B _08424_/Y VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout719 VGND VPWR _12195_/B1 _12121_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_08800_ VGND VPWR VPWR VGND _15209_/D _08814_/S fanout23/X hold1138/X sky130_fd_sc_hd__mux2_4
X_09780_ VGND VPWR VPWR VGND _14269_/D fanout39/X _09792_/S hold908/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Left_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08731_ VGND VPWR VGND VPWR _15268_/D hold1000/X _08731_/A2 _08730_/X _11296_/A sky130_fd_sc_hd__o211a_1
X_08662_ VPWR VGND VPWR VGND _15292_/Q _08667_/A2 _08662_/X _08662_/B1 _08661_/X _08722_/C1
+ sky130_fd_sc_hd__a221o_1
X_07613_ _07614_/C _07609_/X _07611_/X _07612_/Y _07974_/B1 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_08593_ _08995_/B _07494_/X _08604_/B2 _08592_/Y _08591_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07544_ VPWR VGND _07544_/X _07544_/B _15560_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07475_ VGND VPWR VPWR VGND _07479_/A _07703_/A _09164_/A _15591_/Q sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_46_Left_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09214_ VGND VPWR VPWR VGND _14879_/D hold1083/X _09229_/S fanout37/X sky130_fd_sc_hd__mux2_1
X_09145_ VGND VPWR VPWR VGND _14953_/D fanout38/X _09160_/S hold808/X sky130_fd_sc_hd__mux2_1
X_09076_ VGND VPWR VPWR VGND _15017_/D hold979/X _09088_/S fanout38/X sky130_fd_sc_hd__mux2_1
X_14079__1196 VPWR VGND VPWR VGND _15498_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_08027_ VGND VPWR VPWR VGND _08027_/X _10064_/B _08182_/S _12799_/B sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_55_Left_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold762 hold762/X hold762/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 hold740/X hold740/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 hold751/X hold751/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 hold773/X hold773/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 hold795/X hold795/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 hold784/X hold784/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ VPWR VGND VGND VPWR _09967_/Y _12878_/C _09977_/Y _09966_/X _14804_/D sky130_fd_sc_hd__o22ai_1
X_08929_ VPWR VGND VPWR VGND _14150_/Q hold226/A _14151_/Q _09885_/C sky130_fd_sc_hd__or3_1
X_11940_ VGND VPWR VGND VPWR _11940_/X _14485_/Q _12192_/A2 _11948_/S _11939_/X sky130_fd_sc_hd__o211a_1
Xhold1440 _08428_/A _15362_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 hold1451/X hold977/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13199__316 VPWR VGND VPWR VGND _14474_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_79_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1462 hold1462/X _15268_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11871_ VGND VPWR VGND VPWR _11871_/X _11870_/X _11869_/X _12174_/S _12184_/C1 sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_64_Left_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_60_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_55_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14590_ hold207/A _14590_/CLK _14590_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10822_ VGND VPWR VGND VPWR _14398_/D _12602_/B1 _10820_/X _10821_/X _12751_/C1 sky130_fd_sc_hd__o211a_1
X_10753_ VPWR VGND VGND VPWR _10753_/X _11092_/S _10753_/B sky130_fd_sc_hd__or2_1
XFILLER_38_1033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_41_864 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_71_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10684_ VGND VPWR VPWR VGND _10684_/X hold694/A _10687_/B hold242/A sky130_fd_sc_hd__mux2_1
X_15211_ hold230/A _15211_/CLK _15211_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12423_ VPWR VGND VGND VPWR _12423_/X _12655_/S _12423_/B sky130_fd_sc_hd__or2_1
X_12354_ VGND VPWR VPWR VGND _12354_/X _14464_/Q _12370_/S _14752_/Q sky130_fd_sc_hd__mux2_1
X_15142_ _15142_/Q _15142_/CLK _15142_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_73_Left_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11305_ VPWR VGND VGND VPWR _11305_/X _14820_/Q _11307_/B sky130_fd_sc_hd__or2_1
X_15073_ _15073_/Q clkload14/A _15073_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12285_ VGND VPWR VPWR VGND _12285_/X _12282_/X _12684_/S _12281_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_798 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11236_ VGND VPWR VPWR VGND _11236_/X _11233_/X _11244_/S _11232_/X sky130_fd_sc_hd__mux2_1
X_11167_ VGND VPWR VPWR VGND _11167_/X hold656/A _11167_/S hold299/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10118_ VPWR VGND VPWR VGND _10117_/X _10618_/A _12121_/B1 _10118_/X sky130_fd_sc_hd__a21o_1
XFILLER_23_1302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11098_ VGND VPWR VPWR VGND _11098_/X _14438_/Q _11098_/S hold570/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14926_ _14926_/Q clkload28/A _14926_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10049_ VPWR VGND VGND VPWR _10050_/B _15636_/Q _10049_/B sky130_fd_sc_hd__or2_1
XFILLER_36_636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14857_ _14857_/Q clkload28/A _14857_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14788_ hold706/A _14788_/CLK _14788_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_371 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_34_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07260_ VPWR VGND VGND VPWR _07272_/D _08047_/A _07260_/B sky130_fd_sc_hd__nand2_1
X_07191_ VGND VPWR VPWR VGND _07355_/B _11535_/A _07230_/S _14389_/Q sky130_fd_sc_hd__mux2_1
X_15409_ hold650/A _15409_/CLK _15409_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09901_ VPWR VGND VPWR VGND _09893_/Y hold714/X _09907_/S hold715/A _09900_/Y sky130_fd_sc_hd__a22o_1
Xfanout505 VGND VPWR _07568_/X _12227_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout538 VGND VPWR fanout539/X fanout538/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout516 VPWR VGND _12372_/S fanout539/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout527 VGND VPWR fanout538/X _12747_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09832_ VGND VPWR VPWR VGND _14220_/D fanout98/X _09833_/S hold548/X sky130_fd_sc_hd__mux2_1
Xfanout549 VPWR VGND VGND VPWR clone13/A _07558_/B sky130_fd_sc_hd__buf_12
X_09763_ VGND VPWR VPWR VGND _14283_/D fanout97/X _09763_/S hold563/X sky130_fd_sc_hd__mux2_1
X_13690__807 VPWR VGND VPWR VGND _15030_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_08714_ VPWR VGND VPWR VGND hold895/A _08714_/A2 _08714_/X _08664_/X _08665_/X _08726_/C1
+ sky130_fd_sc_hd__a221o_1
X_09694_ VPWR VGND VGND VPWR _09694_/B _09694_/Y _09694_/A sky130_fd_sc_hd__nor2_2
Xrebuffer21 VPWR VGND VPWR VGND _07328_/B _07703_/A sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer10 VPWR VGND VPWR VGND _07144_/A1 _07143_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer32 VPWR VGND VPWR VGND rebuffer32/X rebuffer33/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer43 VPWR VGND VPWR VGND rebuffer43/X _07703_/A sky130_fd_sc_hd__dlygate4sd1_1
X_08645_ VPWR VGND VGND VPWR _08645_/X _14391_/Q _08664_/B sky130_fd_sc_hd__or2_1
X_13911__1028 VPWR VGND VPWR VGND _15283_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_13731__848 VPWR VGND VPWR VGND _15103_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_08576_ VPWR VGND VPWR VGND _08575_/Y _10060_/C _08571_/Y _08986_/B _07534_/B sky130_fd_sc_hd__a22o_1
X_07527_ VPWR VGND _07527_/X _07544_/B _15562_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_23_831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_74_1299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07458_ VPWR VGND VGND VPWR _15452_/Q _15597_/Q _07492_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13584__701 VPWR VGND VPWR VGND _14915_/CLK clkload48/A sky130_fd_sc_hd__inv_2
X_07389_ VPWR VGND VGND VPWR _07389_/A _07389_/Y _07389_/B sky130_fd_sc_hd__nand2_1
X_09128_ VGND VPWR VPWR VGND _14967_/D hold532/X _09128_/S fanout96/X sky130_fd_sc_hd__mux2_1
X_13625__742 VPWR VGND VPWR VGND _14965_/CLK clkload54/A sky130_fd_sc_hd__inv_2
XFILLER_2_724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09059_ VGND VPWR VPWR VGND _15031_/D hold892/X _09059_/S fanout96/X sky130_fd_sc_hd__mux2_1
Xhold570 hold570/X hold570/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 hold581/X hold581/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12070_ VPWR VGND VGND VPWR _12070_/X hold298/A _12219_/S sky130_fd_sc_hd__or2_1
X_12931__48 VPWR VGND VPWR VGND _14174_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_11021_ VGND VPWR VGND VPWR _11021_/X _11185_/A1 _11017_/X _11020_/X _11180_/C1 sky130_fd_sc_hd__o211a_1
Xhold592 hold592/X hold592/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_58_761 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_45_400 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1270 hold1270/X _14561_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1292 hold1292/X _14824_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1281 hold1281/X _15635_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14711_ hold502/A _14711_/CLK _14711_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11923_ VGND VPWR VPWR VGND _11923_/X hold885/A _12149_/S hold836/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11854_ VPWR VGND VGND VPWR _11854_/X hold524/A _12183_/S sky130_fd_sc_hd__or2_1
XFILLER_33_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14642_ hold350/A _14642_/CLK _14642_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10805_ VPWR VGND VPWR VGND _10802_/X _11215_/C1 _10804_/X _10805_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_499 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14573_ hold200/A _14573_/CLK _14573_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11785_ VGND VPWR VGND VPWR _11785_/X _15004_/Q _12188_/A2 _11995_/S _11784_/X sky130_fd_sc_hd__o211a_1
X_10736_ VGND VPWR VGND VPWR _10736_/X _10735_/X _10734_/X _10732_/S _10741_/C1 sky130_fd_sc_hd__a211o_1
X_10667_ VGND VPWR VGND VPWR _10667_/X _10664_/X _10666_/X _10557_/A _10667_/C1 sky130_fd_sc_hd__a211o_1
X_12406_ VGND VPWR VGND VPWR _12406_/X _12405_/X _12404_/X _12721_/S _12720_/C1 sky130_fd_sc_hd__a211o_1
X_15125_ _15125_/Q _15125_/CLK _15125_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10598_ VPWR VGND _10598_/X _10597_/X _10593_/X clone2/A _10589_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12337_ VGND VPWR VGND VPWR _12337_/X _12334_/X _12336_/X _12588_/A1 _12748_/C1 sky130_fd_sc_hd__a211o_1
X_13368__485 VPWR VGND VPWR VGND _14643_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
XFILLER_64_1424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12268_ VPWR VGND VGND VPWR _12249_/X _12266_/X _07913_/Y _12267_/X _12268_/X sky130_fd_sc_hd__o22a_1
X_15056_ hold527/A _15056_/CLK _15056_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11219_ VGND VPWR VPWR VGND _11219_/X _15396_/Q _11223_/S hold325/A sky130_fd_sc_hd__mux2_1
X_12199_ VGND VPWR VPWR VGND _12199_/X hold682/A _12228_/B hold258/A sky130_fd_sc_hd__mux2_1
XFILLER_7_1340 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14909_ hold576/A _14909_/CLK _14909_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_64_786 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08430_ VPWR VGND VGND VPWR _08430_/X hold728/X _08484_/B sky130_fd_sc_hd__or2_1
XFILLER_52_937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14078__1195 VPWR VGND VPWR VGND _15497_/CLK clkload20/A sky130_fd_sc_hd__inv_2
XFILLER_36_488 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_24_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08361_ VGND VPWR VPWR VGND _15412_/D hold488/X _08375_/S fanout26/X sky130_fd_sc_hd__mux2_1
X_07312_ VPWR VGND VGND VPWR _07313_/B _07310_/Y _07812_/A _07813_/A _07859_/A _07820_/A
+ sky130_fd_sc_hd__o41a_1
X_08292_ VPWR VGND VPWR VGND _10061_/D _07574_/A _08291_/X _08292_/X sky130_fd_sc_hd__a21o_1
X_07243_ VPWR VGND _07243_/X _07358_/B _07244_/A _15453_/Q _07241_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_34_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13609__726 VPWR VGND VPWR VGND _14949_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_07174_ VPWR VGND VPWR VGND _07174_/Y _07314_/B sky130_fd_sc_hd__inv_2
Xfanout302 VGND VPWR _10479_/S _10702_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout313 VPWR VGND _10742_/S fanout314/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout324 VGND VPWR _11102_/S _10885_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout346 VGND VPWR _11093_/S _10835_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09815_ VGND VPWR VPWR VGND _14237_/D fanout40/X _09830_/S hold505/X sky130_fd_sc_hd__mux2_1
XFILLER_59_525 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout357 VGND VPWR _10677_/S _10467_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout335 VGND VPWR _11068_/S _11054_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout379 VGND VPWR _11205_/A _11092_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout368 VGND VPWR fanout382/X _11244_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13161__278 VPWR VGND VPWR VGND _14436_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_09746_ VGND VPWR VPWR VGND _14300_/D fanout35/X _09756_/S hold408/X sky130_fd_sc_hd__mux2_1
X_09677_ VGND VPWR VPWR VGND _14363_/D hold1042/X _09684_/S fanout33/X sky130_fd_sc_hd__mux2_1
XFILLER_36_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_76_1317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08628_ VGND VPWR VGND VPWR _15300_/D hold960/X _08628_/A2 _08627_/X _09977_/A sky130_fd_sc_hd__o211a_1
XFILLER_55_775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_43_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08559_ VPWR VGND VGND VPWR _08559_/A _08559_/Y _08559_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11570_ VGND VPWR VPWR VGND _11570_/X hold602/A _12094_/S hold160/A sky130_fd_sc_hd__mux2_1
X_10521_ VPWR VGND VGND VPWR _10521_/X hold343/A _10521_/B sky130_fd_sc_hd__or2_1
X_13055__172 VPWR VGND VPWR VGND _14298_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_10452_ VGND VPWR VGND VPWR _14388_/D _11973_/B _10450_/X _10451_/X _11937_/C1 sky130_fd_sc_hd__o211a_1
X_10383_ VPWR VGND VGND VPWR _10383_/X _10685_/S _10383_/B sky130_fd_sc_hd__or2_1
X_12122_ VPWR VGND VGND VPWR _12103_/Y _12121_/X _10710_/B _15459_/Q _15459_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
X_12053_ VPWR VGND VGND VPWR _12053_/X _12069_/S _12053_/B sky130_fd_sc_hd__or2_1
XFILLER_77_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11004_ VGND VPWR VGND VPWR _11004_/X _11001_/X _11003_/X _11004_/A1 _11237_/A1 sky130_fd_sc_hd__a211o_1
X_13402__519 VPWR VGND VPWR VGND _14677_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_46_1198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout880 VPWR VGND _09164_/A _15578_/Q VPWR VGND sky130_fd_sc_hd__buf_2
Xclkbuf_3_6_0_clk clkload4/A clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_24_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13753__870 VPWR VGND VPWR VGND _15125_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11906_ VGND VPWR VGND VPWR _11906_/X _12156_/A1 _11902_/X _11905_/X _12202_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_34_948 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11837_ VGND VPWR VPWR VGND _11837_/X _14194_/Q _11838_/S hold225/A sky130_fd_sc_hd__mux2_1
X_14625_ _14625_/Q _14625_/CLK _14625_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_42_981 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14556_ hold584/A _14556_/CLK _14556_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11768_ VPWR VGND VPWR VGND _11767_/X _12101_/A1 _11766_/X _11768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10719_ VPWR VGND VPWR VGND _10718_/X _10745_/C1 _10717_/X _10719_/Y sky130_fd_sc_hd__a21oi_1
X_14487_ hold763/A _14487_/CLK _14487_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11699_ VGND VPWR VPWR VGND _11699_/X _11698_/X _12476_/S _11697_/X sky130_fd_sc_hd__mux2_1
Xrebuffer1 rebuffer1/X _07557_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_15108_ _15108_/Q _15108_/CLK _15108_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13910__1027 VPWR VGND VPWR VGND _15282_/CLK clkload17/A sky130_fd_sc_hd__inv_2
X_07930_ VPWR VGND VPWR VGND _07962_/A _15561_/Q _15562_/Q _07931_/B sky130_fd_sc_hd__a21oi_1
X_15039_ hold616/A _15039_/CLK _15039_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07861_ VPWR VGND VPWR VGND _15087_/Q _07881_/A2 _07861_/X _07668_/B _07298_/A _07860_/Y
+ sky130_fd_sc_hd__a221o_1
X_07792_ VPWR VGND VPWR VGND _07730_/B _15558_/Q _07999_/A _07992_/A sky130_fd_sc_hd__a21o_1
X_09600_ VGND VPWR VPWR VGND _14468_/D fanout66/X _09619_/S hold587/X sky130_fd_sc_hd__mux2_1
XFILLER_49_591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09531_ VGND VPWR VPWR VGND _14531_/D fanout63/X _09552_/S hold179/X sky130_fd_sc_hd__mux2_1
X_09462_ VGND VPWR VPWR VGND _14594_/D fanout58/X _09467_/S hold336/X sky130_fd_sc_hd__mux2_1
X_08413_ VPWR VGND VGND VPWR _14810_/Q hold153/A _08413_/Y sky130_fd_sc_hd__nor2_1
X_09393_ VGND VPWR VPWR VGND _14656_/D hold379/X _09411_/S fanout48/X sky130_fd_sc_hd__mux2_1
XFILLER_36_1312 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_52_789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08344_ _15429_/D fanout92/X fanout88/X _08356_/S _08343_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_13039__156 VPWR VGND VPWR VGND _14282_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_08275_ VPWR VGND _08275_/X _08275_/B _08275_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_07226_ VPWR VGND VPWR VGND _07226_/Y _07360_/A _07224_/X _07110_/Y _07143_/X sky130_fd_sc_hd__a211oi_1
X_07157_ VPWR VGND VGND VPWR _15474_/Q _07157_/B _07626_/A sky130_fd_sc_hd__nor2_1
X_07088_ VPWR VGND VPWR VGND _07088_/Y _15458_/Q sky130_fd_sc_hd__inv_2
X_13696__813 VPWR VGND VPWR VGND _15036_/CLK clkload11/A sky130_fd_sc_hd__inv_2
Xfanout110 VGND VPWR _09726_/A1 _08266_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout121 VPWR VGND _09862_/A0 _09723_/A1 VPWR VGND sky130_fd_sc_hd__buf_4
X_12901__18 VPWR VGND VPWR VGND _14143_/CLK clkload29/A sky130_fd_sc_hd__inv_2
Xfanout154 VPWR VGND _08969_/A _08972_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout132 VPWR VGND VGND VPWR clone17/A _07914_/B1 sky130_fd_sc_hd__buf_8
Xfanout143 VPWR VGND _08721_/A2 _08704_/A2 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout165 VGND VPWR _11625_/S _12100_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_75_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13737__854 VPWR VGND VPWR VGND _15109_/CLK clkload46/A sky130_fd_sc_hd__inv_2
XFILLER_47_517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xfanout198 VGND VPWR _11638_/A1 _12119_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout187 VGND VPWR _12536_/S _12665_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout176 VGND VPWR _12069_/S _12221_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09729_ VPWR VGND VGND VPWR _09799_/B _09729_/Y _09729_/A sky130_fd_sc_hd__nor2_2
XFILLER_76_1103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_femto_892 uio_oe[3] tt_um_femto_892/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_12740_ VGND VPWR VGND VPWR _12740_/X _12740_/A1 _12735_/X _12739_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_12671_ VGND VPWR VPWR VGND _12671_/X hold510/A _12671_/S hold624/A sky130_fd_sc_hd__mux2_1
XFILLER_70_597 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_63_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14410_ _14410_/Q clkload33/A _14410_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11622_ VPWR VGND VGND VPWR _12103_/A _11622_/B _11622_/Y sky130_fd_sc_hd__nor2_1
X_15390_ hold810/A _15390_/CLK _15390_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14341_ hold946/A _14341_/CLK _14341_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11553_ VGND VPWR _11551_/B _15437_/Q _11553_/Y _11551_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_10_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14272_ hold999/A _14272_/CLK _14272_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11484_ VGND VPWR VPWR VGND _11484_/X _15080_/Q _11490_/S _15078_/Q sky130_fd_sc_hd__mux2_1
X_10504_ VGND VPWR VPWR VGND _10504_/X _10501_/X _10510_/S _10500_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_668 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10435_ VPWR VGND VPWR VGND _10432_/X _10557_/A _10434_/X _10435_/X sky130_fd_sc_hd__a21o_1
X_14077__1194 VPWR VGND VPWR VGND _15496_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_10366_ VGND VPWR VGND VPWR _10366_/X _10365_/X _10364_/X _10615_/S _10622_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_3_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12105_ VGND VPWR VPWR VGND _12105_/X hold949/A _12117_/B hold724/A sky130_fd_sc_hd__mux2_1
X_10297_ VGND VPWR VGND VPWR _10297_/X _10294_/X _10296_/X _10523_/A1 _10634_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_66_804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12036_ VGND VPWR VGND VPWR _12036_/X _12035_/X _12034_/X _12118_/B1 _12115_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_61_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_59_1345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_61_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12869_ VGND VPWR VPWR VGND _15593_/D _12869_/A1 _12870_/S _15593_/Q sky130_fd_sc_hd__mux2_1
X_14608_ hold784/A _14608_/CLK _14608_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13530__647 VPWR VGND VPWR VGND _14810_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_15588_ _15588_/Q clkload44/A _15588_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14539_ hold803/A _14539_/CLK _14539_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08060_ VPWR VGND VGND VPWR _08220_/A _08060_/B _08060_/Y sky130_fd_sc_hd__nor2_1
X_12967__84 VPWR VGND VPWR VGND _14210_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_13383__500 VPWR VGND VPWR VGND _14658_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_08962_ VGND VPWR VPWR VGND _08963_/B _07533_/X _09906_/A hold888/A sky130_fd_sc_hd__mux2_1
X_13424__541 VPWR VGND VPWR VGND _14699_/CLK clkload12/A sky130_fd_sc_hd__inv_2
X_08893_ VGND VPWR VGND VPWR _15146_/D hold1411/X _08893_/A2 _08892_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_07913_ VPWR VGND VPWR VGND _07913_/Y _12584_/A sky130_fd_sc_hd__inv_4
X_07844_ VGND VPWR _07864_/A _15564_/Q _15565_/Q _07906_/A VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_77_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07775_ VPWR VGND VPWR VGND _08218_/B _07761_/B _07759_/X _08210_/A sky130_fd_sc_hd__a21o_1
Xclone6 VGND VPWR clone6/A clone6/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09514_ VGND VPWR VPWR VGND _14545_/D _09827_/A1 _09514_/S hold1013/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09445_ VGND VPWR VPWR VGND _14607_/D _09863_/A0 _09446_/S hold746/X sky130_fd_sc_hd__mux2_1
XFILLER_24_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09376_ VGND VPWR VPWR VGND _14670_/D hold672/X _09376_/S _09690_/A0 sky130_fd_sc_hd__mux2_1
X_08327_ VGND VPWR VPWR VGND _15492_/D _08091_/X _08338_/S hold669/X sky130_fd_sc_hd__mux2_1
X_08258_ VGND VPWR _08258_/X _08258_/B _10061_/A _08275_/A VPWR VGND sky130_fd_sc_hd__and3_1
X_07209_ VPWR VGND _07209_/X _07372_/C _15451_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_08189_ VGND VPWR _08188_/X _10059_/A _08189_/Y _08185_/Y VPWR VGND sky130_fd_sc_hd__o21ai_2
X_10220_ VGND VPWR VPWR VGND _10220_/X hold719/A _11231_/S hold290/A sky130_fd_sc_hd__mux2_1
XFILLER_0_822 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10151_ VPWR VGND VGND VPWR _10151_/X hold549/A _10604_/S sky130_fd_sc_hd__or2_1
XFILLER_58_55 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10082_ VPWR VGND _14153_/D _11340_/A _10081_/Y _10056_/A _10079_/X _10080_/X VPWR
+ VGND sky130_fd_sc_hd__a311oi_1
X_13167__284 VPWR VGND VPWR VGND _14442_/CLK clkload33/A sky130_fd_sc_hd__inv_2
X_14890_ _14890_/Q _14890_/CLK _14890_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_63_807 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10984_ VGND VPWR VGND VPWR _10984_/X _11004_/A1 _10980_/X _10983_/X _11235_/C1 sky130_fd_sc_hd__o211a_1
X_15511_ hold814/A _15511_/CLK _15511_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12723_ VGND VPWR VPWR VGND _12727_/B _14799_/Q _12736_/B _14250_/Q sky130_fd_sc_hd__mux2_1
XFILLER_43_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15442_ _15442_/Q clkload47/A _15442_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12654_ VGND VPWR VGND VPWR _12654_/X _12662_/A1 _12650_/X _12653_/X _12662_/C1 sky130_fd_sc_hd__o211a_1
X_12585_ VPWR VGND VGND VPWR _12585_/X _15425_/Q _12599_/S sky130_fd_sc_hd__or2_1
X_15373_ hold486/A _15373_/CLK _15373_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1395 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11605_ VGND VPWR VPWR VGND _11609_/B hold519/A _12097_/S hold460/A sky130_fd_sc_hd__mux2_1
X_13865__982 VPWR VGND VPWR VGND _15237_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_11536_ VPWR VGND _11536_/X _10072_/B _15095_/Q _10072_/A _11535_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14324_ hold773/A _14324_/CLK _14324_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14255_ hold703/A _14255_/CLK _14255_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11467_ VGND VPWR VPWR VGND _11467_/X _11466_/X _11476_/S _15453_/Q sky130_fd_sc_hd__mux2_1
X_11398_ _11400_/A _14851_/Q _11398_/A _14852_/Q _11398_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_14186_ _14186_/Q _14186_/CLK _14186_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13408__525 VPWR VGND VPWR VGND _14683_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_10418_ VGND VPWR VPWR VGND _10418_/X _10417_/X _10652_/S _10416_/X sky130_fd_sc_hd__mux2_1
X_14809__937 _14809_/D _14809__937/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_10349_ VPWR VGND VPWR VGND _10348_/X _10608_/A1 _10347_/X _10349_/Y sky130_fd_sc_hd__a21oi_1
X_12019_ VPWR VGND VPWR VGND _12018_/X _12193_/C1 _12017_/X _12019_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_1344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_66_634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07560_ VGND VPWR VGND VPWR _07559_/A _07560_/X _07560_/D _07560_/C _07560_/B sky130_fd_sc_hd__and4b_4
XFILLER_53_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_62_840 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1059 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07491_ _07492_/B _07489_/B _07489_/A _08603_/A _07462_/A _08597_/A VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__o311a_1
X_09230_ VGND VPWR VPWR VGND _14863_/D hold1136/X _09231_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
X_09161_ VGND VPWR VPWR VGND _14937_/D _09229_/A0 _09161_/S hold948/X sky130_fd_sc_hd__mux2_1
XFILLER_72_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08112_ VPWR VGND VPWR VGND _08112_/Y _08112_/A sky130_fd_sc_hd__inv_2
X_09092_ VGND VPWR VPWR VGND _15001_/D hold1022/X _09092_/S _09229_/A0 sky130_fd_sc_hd__mux2_1
X_08043_ VGND VPWR VGND VPWR _07380_/X _07254_/Y _08064_/B _08044_/B sky130_fd_sc_hd__o21ba_1
Xhold911 hold911/X hold911/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold900 hold900/X hold900/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 hold922/X hold922/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 hold944/X hold944/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 hold933/X hold933/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 hold955/X hold955/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 hold988/X hold988/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ VPWR VGND VGND VPWR _09996_/C _09994_/B _15612_/D sky130_fd_sc_hd__nor2_1
Xhold977 hold977/X hold977/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 hold966/X hold966/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 hold999/X hold999/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08945_ VPWR VGND _15125_/D _08945_/B _08955_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_69_472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08876_ VPWR VGND VGND VPWR _08876_/X _15154_/Q _08926_/B sky130_fd_sc_hd__or2_1
X_07827_ VGND VPWR VPWR VGND _07827_/D _07827_/C _07827_/B _07827_/A _12831_/A sky130_fd_sc_hd__or4_4
X_13201__318 VPWR VGND VPWR VGND _14476_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_07758_ VPWR VGND VPWR VGND _07826_/D _15594_/Q _10078_/A _07760_/B _09240_/A sky130_fd_sc_hd__a22o_1
X_14076__1193 VPWR VGND VPWR VGND _15495_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_07689_ VGND VPWR VPWR VGND _15538_/D fanout67/X _08231_/S hold272/X sky130_fd_sc_hd__mux2_1
X_09428_ VGND VPWR VPWR VGND _09446_/S fanout48/X hold1202/X _14624_/D sky130_fd_sc_hd__mux2_2
X_13849__966 VPWR VGND VPWR VGND _15221_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_09359_ VGND VPWR VPWR VGND _14687_/D hold565/X _09376_/S fanout45/X sky130_fd_sc_hd__mux2_1
XFILLER_40_556 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12370_ VGND VPWR VPWR VGND _12370_/X _15020_/Q _12370_/S hold748/A sky130_fd_sc_hd__mux2_1
X_11321_ VPWR VGND VGND VPWR _11342_/C _14826_/Q _14825_/Q sky130_fd_sc_hd__or2_1
X_11252_ VGND VPWR VGND VPWR _11252_/X _14966_/Q _11252_/A2 _11251_/X _11252_/C1 sky130_fd_sc_hd__o211a_1
X_10203_ VGND VPWR VPWR VGND _10203_/X hold492/A _10567_/S hold259/A sky130_fd_sc_hd__mux2_1
X_11183_ VPWR VGND VGND VPWR _11183_/X hold208/A _11186_/S sky130_fd_sc_hd__or2_1
X_10134_ VGND VPWR VPWR VGND _10134_/X _10131_/X _10615_/S _10130_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10065_ _10064_/X _10065_/B _10065_/X _10065_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_14942_ _14942_/Q _14942_/CLK _14942_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1006 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14873_ hold994/A _14873_/CLK _14873_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10967_ VGND VPWR VGND VPWR _10967_/X _10964_/X _10966_/X _11189_/A1 _11245_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_43_372 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12706_ VGND VPWR VPWR VGND _12706_/X hold814/A _12708_/S hold210/A sky130_fd_sc_hd__mux2_1
XFILLER_31_545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10898_ VGND VPWR VPWR VGND _10898_/X _14497_/Q _10919_/S hold628/A sky130_fd_sc_hd__mux2_1
X_15425_ _15425_/Q _15425_/CLK _15425_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12637_ VGND VPWR VGND VPWR _12637_/X _12634_/X _12636_/X _12624_/S _12739_/C1 sky130_fd_sc_hd__a211o_1
X_12568_ VGND VPWR VPWR VGND _12568_/X _14502_/Q _12578_/S _14182_/Q sky130_fd_sc_hd__mux2_1
X_15356_ _15356_/Q _15356_/CLK _15356_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold207 hold207/X hold207/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_15287_ hold952/A _15287_/CLK _15287_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12937__54 VPWR VGND VPWR VGND _14180_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_11519_ VGND VPWR VPWR VGND _15090_/D _11518_/X _11528_/S _15090_/Q sky130_fd_sc_hd__mux2_1
X_12499_ VGND VPWR VPWR VGND _12499_/X _12496_/X _12665_/S _12495_/X sky130_fd_sc_hd__mux2_1
X_14307_ hold293/A _14307_/CLK _14307_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14238_ hold268/A _14238_/CLK _14238_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold218 hold218/X hold218/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold229/X hold229/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14169_ hold351/A _14169_/CLK _14169_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13642__759 VPWR VGND VPWR VGND _14982_/CLK clkload17/A sky130_fd_sc_hd__inv_2
Xfanout709 VGND VPWR _08484_/B _08482_/B VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_13495__612 VPWR VGND VPWR VGND _14770_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_08730_ VGND VPWR VGND VPWR _08730_/X _08522_/B _08730_/B1 _14379_/Q _08523_/B sky130_fd_sc_hd__a211o_1
X_08661_ VPWR VGND VGND VPWR _08660_/X _08690_/S _08194_/Y _14404_/Q _08661_/X _08659_/Y
+ sky130_fd_sc_hd__o221a_1
X_07612_ VPWR VGND VGND VPWR _07612_/A _10075_/A _07612_/Y sky130_fd_sc_hd__nor2_1
X_08592_ VPWR VGND VGND VPWR _08592_/A _08592_/B _08592_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13536__653 VPWR VGND VPWR VGND _14867_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_07543_ VGND VPWR VGND VPWR _07542_/X _08956_/B _07534_/B _15564_/Q _07541_/Y _08943_/A
+ sky130_fd_sc_hd__o221ai_4
X_07474_ VPWR VGND VGND VPWR _15447_/Q _07483_/A _07482_/B sky130_fd_sc_hd__nand2_1
X_09213_ VGND VPWR VPWR VGND _14880_/D hold868/X _09213_/S _07953_/X sky130_fd_sc_hd__mux2_1
X_09144_ VGND VPWR VPWR VGND _14954_/D clone6/A _09160_/S hold743/X sky130_fd_sc_hd__mux2_1
X_09075_ VGND VPWR VPWR VGND _15018_/D hold1043/X _09088_/S fanout41/X sky130_fd_sc_hd__mux2_1
X_08026_ VGND VPWR _08026_/B _10064_/B _08026_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold730 hold730/X hold730/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 hold741/X hold741/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 hold763/X hold763/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 hold752/X hold752/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 hold785/X hold785/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 hold774/X hold774/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 hold796/X hold796/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09977_ VPWR VGND VGND VPWR _09977_/A _09977_/Y _09977_/B sky130_fd_sc_hd__nand2_1
X_08928_ VGND VPWR VGND VPWR _08935_/A clone20/A _15638_/Q _15479_/Q sky130_fd_sc_hd__a21bo_1
XFILLER_57_431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1430 hold1430/X _14186_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 hold1452/X hold883/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 hold1441/X _15281_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08859_ VGND VPWR VPWR VGND hold714/A _08859_/C _14144_/Q _09900_/A sky130_fd_sc_hd__or3_2
Xhold1463 _08872_/A _15156_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11870_ VGND VPWR VPWR VGND _11870_/X hold522/A _12183_/S hold178/A sky130_fd_sc_hd__mux2_1
X_10821_ VPWR VGND VGND VPWR _10821_/X _14398_/Q _12269_/B sky130_fd_sc_hd__or2_1
XFILLER_38_1023 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13279__396 VPWR VGND VPWR VGND _14554_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_10752_ VGND VPWR VPWR VGND _10752_/X hold479/A _10835_/B hold256/A sky130_fd_sc_hd__mux2_1
XFILLER_9_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10683_ VGND VPWR VPWR VGND _10683_/X _14203_/Q _10687_/B hold230/A sky130_fd_sc_hd__mux2_1
X_15210_ hold328/A _15210_/CLK _15210_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12422_ VGND VPWR VPWR VGND _12422_/X hold603/A _12661_/S hold336/A sky130_fd_sc_hd__mux2_1
X_12353_ VGND VPWR VPWR VGND _12353_/X _14208_/Q _12370_/S _15216_/Q sky130_fd_sc_hd__mux2_1
X_15141_ _15141_/Q _15141_/CLK _15141_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11304_ VGND VPWR VGND VPWR _14819_/D _14379_/Q _11303_/B _11303_/Y _11315_/A1 sky130_fd_sc_hd__o211a_1
X_12284_ VGND VPWR VGND VPWR _12284_/X _12256_/S _12280_/X _12283_/X _12702_/C1 sky130_fd_sc_hd__o211a_1
X_15072_ _15072_/Q clkload15/A _15072_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11235_ VGND VPWR VGND VPWR _11235_/X _11235_/A1 _11231_/X _11234_/X _11235_/C1 sky130_fd_sc_hd__o211a_1
X_11166_ VGND VPWR VPWR VGND _11166_/X _14216_/Q _11167_/S hold171/A sky130_fd_sc_hd__mux2_1
X_11097_ VGND VPWR VGND VPWR _11097_/X _11104_/B1 _11092_/X _11096_/X _10765_/S sky130_fd_sc_hd__o211a_1
X_10117_ VPWR VGND _10117_/X _10116_/X _10112_/X _10617_/S _10108_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_10048_ VPWR VGND VGND VPWR _15636_/Q _10051_/B _10049_/B sky130_fd_sc_hd__nand2_1
X_14925_ _14925_/Q _14925_/CLK _14925_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13223__340 VPWR VGND VPWR VGND _14498_/CLK clkload42/A sky130_fd_sc_hd__inv_2
XFILLER_76_784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14856_ _14856_/Q clkload28/A _14856_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14787_ hold438/A _14787_/CLK _14787_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_51_629 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11999_ VGND VPWR VGND VPWR _11999_/X _11998_/X _11997_/X _11995_/S _12017_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_16_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15408_ hold699/A _15408_/CLK _15408_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07190_ VGND VPWR VGND VPWR _07188_/X _08083_/A _07190_/B sky130_fd_sc_hd__nand2b_2
X_15339_ _15339_/Q _15339_/CLK _15339_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13072__189 VPWR VGND VPWR VGND _14315_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XFILLER_8_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09900_ VPWR VGND VGND VPWR _09900_/A _09900_/Y _09900_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout506 VGND VPWR _12477_/B _12052_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_14075__1192 VPWR VGND VPWR VGND _15494_/CLK clkload16/A sky130_fd_sc_hd__inv_2
Xfanout539 VGND VPWR _07568_/X fanout539/X VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09831_ VGND VPWR VPWR VGND _14221_/D _09865_/A0 _09833_/S hold257/X sky130_fd_sc_hd__mux2_1
Xfanout528 VGND VPWR fanout538/X _12708_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout517 VGND VPWR _12635_/B _12623_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_80_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09762_ VGND VPWR VPWR VGND _14284_/D fanout99/X _09763_/S hold541/X sky130_fd_sc_hd__mux2_1
XFILLER_41_1414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08713_ VGND VPWR VGND VPWR _15277_/D hold872/X _08721_/A2 _08712_/X _08717_/C1 sky130_fd_sc_hd__o211a_1
Xrebuffer11 VPWR VGND VPWR VGND _07469_/S _07477_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_09693_ VGND VPWR VPWR VGND _14347_/D hold851/X _09693_/S _08299_/X sky130_fd_sc_hd__mux2_1
Xrebuffer33 VPWR VGND VPWR VGND rebuffer33/X rebuffer34/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_445 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xrebuffer22 VPWR VGND VPWR VGND _07563_/A rebuffer23/X sky130_fd_sc_hd__dlygate4sd1_1
X_08644_ VGND VPWR VGND VPWR _08714_/A2 _14383_/Q _08194_/B _08644_/X sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_16_Left_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08575_ VGND VPWR _08575_/B _08575_/Y _08575_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_13770__887 VPWR VGND VPWR VGND _15142_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_07526_ VPWR VGND VGND VPWR _07526_/A _07526_/B _07555_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_1332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_640 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07457_ VPWR VGND VGND VPWR _15452_/Q _08597_/A _15597_/Q sky130_fd_sc_hd__nand2_1
X_07388_ VPWR VGND _07397_/A _07899_/B _07389_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_09127_ VGND VPWR VPWR VGND _14968_/D hold549/X _09128_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
X_09058_ VGND VPWR VPWR VGND _15032_/D hold727/X _09059_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
X_13664__781 VPWR VGND VPWR VGND _15004_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_08009_ VGND VPWR VGND VPWR _08009_/X _08005_/Y _08008_/X _08240_/A _07333_/Y sky130_fd_sc_hd__a211o_1
Xhold571 hold571/X hold571/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 hold560/X hold560/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ VPWR VGND VGND VPWR _11020_/X _11176_/S _11020_/B sky130_fd_sc_hd__or2_1
Xhold582 hold582/X hold582/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 hold593/X hold593/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13207__324 VPWR VGND VPWR VGND _14482_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
XFILLER_79_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1260 hold1260/X _14278_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1271 hold1271/X _14342_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 hold1293/X _15146_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 hold1282/X _15362_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14710_ hold870/A _14710_/CLK _14710_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11922_ VGND VPWR VGND VPWR _11922_/X _11921_/X _11920_/X _12156_/A1 _12202_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_79_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14641_ hold606/A _14641_/CLK _14641_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11853_ VGND VPWR VPWR VGND _11853_/X hold562/A _12191_/B hold747/A sky130_fd_sc_hd__mux2_1
X_10804_ VPWR VGND VPWR VGND _10803_/X _11213_/S _11218_/A1 _10804_/X sky130_fd_sc_hd__a21o_1
X_14572_ hold342/A _14572_/CLK _14572_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14099__1216 VPWR VGND VPWR VGND _15518_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_11784_ VPWR VGND VGND VPWR _11784_/X hold433/A _12112_/S sky130_fd_sc_hd__or2_1
X_10735_ VGND VPWR VPWR VGND _10735_/X _14879_/Q _10735_/S hold591/A sky130_fd_sc_hd__mux2_1
X_10666_ VGND VPWR VGND VPWR _10666_/X _15014_/Q _10744_/A2 _10665_/X _10652_/S sky130_fd_sc_hd__o211a_1
X_12405_ VGND VPWR VPWR VGND _12405_/X hold966/A _12409_/B hold590/A sky130_fd_sc_hd__mux2_1
X_15124_ _15124_/Q _15124_/CLK _15124_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10597_ VGND VPWR VGND VPWR _10597_/X _10594_/X _10596_/X _10745_/A1 _10745_/C1 sky130_fd_sc_hd__a211o_1
X_12907__24 VPWR VGND VPWR VGND _14149_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_12336_ VGND VPWR VGND VPWR _12336_/X hold963/A _12705_/A2 _12591_/S _12335_/X sky130_fd_sc_hd__o211a_1
X_12267_ VPWR VGND _12267_/X _12241_/X _12237_/X _12740_/C1 _12584_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_15055_ hold542/A _15055_/CLK _15055_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11218_ VGND VPWR VGND VPWR _11218_/X _11218_/A1 _11213_/X _11217_/X _11218_/C1 sky130_fd_sc_hd__o211a_1
X_12198_ VGND VPWR VPWR VGND _12198_/X hold974/A _12228_/B hold422/A sky130_fd_sc_hd__mux2_1
X_11149_ VGND VPWR VPWR VGND _11149_/X hold537/A _11251_/B hold655/A sky130_fd_sc_hd__mux2_1
X_14908_ hold430/A _14908_/CLK _14908_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14839_ _14839_/Q clkload28/A _14839_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_37_979 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13000__117 VPWR VGND VPWR VGND _14243_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_08360_ VGND VPWR VPWR VGND _15413_/D hold375/X _08375_/S fanout27/X sky130_fd_sc_hd__mux2_1
X_07311_ VPWR VGND VGND VPWR _07311_/A _07311_/B _07812_/A sky130_fd_sc_hd__nor2_1
X_08291_ VPWR VGND VGND VPWR _15445_/Q _08290_/B _08278_/B _08291_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07242_ VPWR VGND VGND VPWR _15454_/Q _07244_/B _07376_/B sky130_fd_sc_hd__nand2_1
X_13648__765 VPWR VGND VPWR VGND _14988_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_07173_ VPWR VGND VGND VPWR _15470_/Q _07173_/B _07314_/B sky130_fd_sc_hd__nor2_1
Xfanout314 VGND VPWR _07893_/X fanout314/X VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout303 VGND VPWR _10479_/S _10700_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout347 VGND VPWR _10795_/S _11093_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout325 VPWR VGND _11102_/S _11241_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_09814_ VGND VPWR VPWR VGND _14238_/D clone6/X _09830_/S hold268/X sky130_fd_sc_hd__mux2_1
Xfanout336 VPWR VGND _11068_/S _10964_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout369 VGND VPWR _10333_/A _11110_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout358 VGND VPWR _10703_/A _10677_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09745_ VGND VPWR VPWR VGND _14301_/D fanout40/X _09757_/S hold183/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_55_721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09676_ VGND VPWR VPWR VGND _14364_/D hold913/X _09684_/S fanout36/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08627_ VPWR VGND VPWR VGND _15299_/Q _08626_/A _08627_/X _08232_/B _08626_/Y _08627_/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_43_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08558_ VGND VPWR VGND VPWR _15314_/D hold942/X _08628_/A2 _08557_/X _11337_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_42_459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08489_ VGND VPWR VGND VPWR _15332_/D input3/X _08458_/B _08488_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
X_07509_ VPWR VGND VGND VPWR _07551_/A _07551_/B _07547_/A _07509_/C sky130_fd_sc_hd__nand3_1
XFILLER_23_673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_1340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10520_ VGND VPWR VPWR VGND _10520_/X hold367/A _10520_/S hold796/A sky130_fd_sc_hd__mux2_1
XFILLER_23_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10451_ VPWR VGND VGND VPWR _10451_/X _14388_/Q _10562_/B sky130_fd_sc_hd__or2_1
XFILLER_10_356 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_1335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10382_ VGND VPWR VPWR VGND _10382_/X hold522/A _10696_/S hold178/A sky130_fd_sc_hd__mux2_1
X_12121_ VPWR VGND VPWR VGND _12120_/X _12029_/A _12121_/B1 _12121_/X sky130_fd_sc_hd__a21o_1
X_14215__933 _14215_/D _14215__933/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_12052_ VGND VPWR VPWR VGND _12052_/X hold640/A _12052_/S hold260/A sky130_fd_sc_hd__mux2_1
Xhold390 hold390/X hold390/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ VGND VPWR VGND VPWR _11003_/X _15023_/Q _11003_/A2 _11002_/X _10985_/S sky130_fd_sc_hd__o211a_1
X_13441__558 VPWR VGND VPWR VGND _14716_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
Xfanout870 VGND VPWR _07511_/B _15601_/Q VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout881 VPWR VGND _12878_/A _15576_/Q VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_24_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1090 hold1090/X _14483_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13294__411 VPWR VGND VPWR VGND _14569_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_11905_ VPWR VGND VGND VPWR _11905_/X _12147_/S _11905_/B sky130_fd_sc_hd__or2_1
XFILLER_61_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14624_ _14624_/Q _14624_/CLK _14624_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11836_ VGND VPWR VPWR VGND _11836_/X hold529/A _12171_/S hold431/A sky130_fd_sc_hd__mux2_1
X_14074__1191 VPWR VGND VPWR VGND _15493_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_14555_ hold613/A _14555_/CLK _14555_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13335__452 VPWR VGND VPWR VGND _14610_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_11767_ VGND VPWR VPWR VGND _11767_/X _11764_/X _12098_/A _11763_/X sky130_fd_sc_hd__mux2_1
X_10718_ VGND VPWR VPWR VGND _10718_/X _10715_/X _10732_/S _10714_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14486_ hold795/A _14486_/CLK _14486_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11698_ VGND VPWR VPWR VGND _11698_/X _14350_/Q _12477_/B hold468/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10649_ VGND VPWR VPWR VGND _10649_/X hold566/A _10670_/S hold193/A sky130_fd_sc_hd__mux2_1
X_15107_ hold920/A _15107_/CLK hold921/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12319_ VGND VPWR VPWR VGND _12319_/X hold573/A _12577_/S hold217/A sky130_fd_sc_hd__mux2_1
X_15038_ hold747/A _15038_/CLK _15038_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07860_ VPWR VGND VGND VPWR _07860_/A _08104_/B _07860_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07791_ VPWR VGND VPWR VGND _07798_/A _07999_/A _07998_/B _07998_/C sky130_fd_sc_hd__a21boi_1
XFILLER_77_890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09530_ VGND VPWR VPWR VGND _14532_/D fanout64/X _09549_/S hold295/X sky130_fd_sc_hd__mux2_1
X_09461_ VGND VPWR VPWR VGND _14595_/D fanout61/X _09482_/S hold269/X sky130_fd_sc_hd__mux2_1
XFILLER_18_990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08412_ VPWR VGND VGND VPWR _14807_/Q _14806_/Q _14808_/Q _09232_/B sky130_fd_sc_hd__o21a_1
XFILLER_52_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09392_ VGND VPWR VPWR VGND _14657_/D hold450/X _09411_/S clone5/X sky130_fd_sc_hd__mux2_1
X_13078__195 VPWR VGND VPWR VGND _14321_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_08343_ VPWR VGND VGND VPWR hold1358/X _08356_/S _08343_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_33_993 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08274_ VPWR VGND VGND VPWR _08290_/A _10061_/B _08275_/B _08290_/B sky130_fd_sc_hd__nand3_1
X_07225_ VPWR VGND VPWR VGND _07143_/X _14380_/Q _07223_/X _07360_/B sky130_fd_sc_hd__a21o_1
X_13882__999 VPWR VGND VPWR VGND _15254_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07156_ VPWR VGND _07159_/A _07157_/B _15474_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07087_ VPWR VGND VPWR VGND _07087_/Y _15465_/Q sky130_fd_sc_hd__inv_2
X_12898__15 VPWR VGND VPWR VGND _14140_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
Xfanout111 VGND VPWR _09229_/A0 _09691_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout100 VGND VPWR _08284_/X _09692_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout122 VPWR VGND _09723_/A1 _08212_/X VPWR VGND sky130_fd_sc_hd__buf_4
X_14098__1215 VPWR VGND VPWR VGND _15517_/CLK clkload35/A sky130_fd_sc_hd__inv_2
Xfanout155 VPWR VGND _08972_/A _08937_/Y VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout133 VPWR VGND clone17/A _07598_/Y VPWR VGND sky130_fd_sc_hd__buf_6
Xfanout144 VGND VPWR _08731_/A2 _08704_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_13776__893 VPWR VGND VPWR VGND _15148_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
Xfanout199 VPWR VGND _11638_/A1 _12226_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout166 VPWR VGND _11625_/S _12118_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout188 VPWR VGND _12536_/S _12373_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout177 VPWR VGND _12069_/S _08298_/A1 VPWR VGND sky130_fd_sc_hd__buf_2
X_07989_ VPWR VGND VPWR VGND _08023_/A _15558_/Q _15559_/Q _07990_/B sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09728_ VGND VPWR VPWR VGND _14315_/D fanout95/X _09728_/S hold602/X sky130_fd_sc_hd__mux2_1
Xtt_um_femto_893 uio_oe[4] tt_um_femto_893/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_76_1115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13319__436 VPWR VGND VPWR VGND _14594_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_09659_ VGND VPWR VPWR VGND _14411_/D hold878/X _09659_/S fanout96/X sky130_fd_sc_hd__mux2_1
XFILLER_63_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_54_1402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12670_ VGND VPWR VGND VPWR _12670_/X _12667_/X _12669_/X _12670_/A1 _12670_/C1 sky130_fd_sc_hd__a211o_1
X_12992__109 VPWR VGND VPWR VGND _14235_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_11621_ VGND VPWR VPWR VGND _11622_/B _11620_/Y _12102_/S _11612_/Y sky130_fd_sc_hd__mux2_1
XFILLER_51_790 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_1419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14340_ hold662/A _14340_/CLK _14340_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11552_ VPWR VGND VPWR VGND _11551_/Y _11274_/B _11542_/A _15436_/D sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14271_ hold970/A _14271_/CLK _14271_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11483_ VGND VPWR VPWR VGND _15078_/D _11482_/X _11492_/S _15078_/Q sky130_fd_sc_hd__mux2_1
X_10503_ VGND VPWR VGND VPWR _10503_/X _10523_/A1 _10499_/X _10502_/X _10630_/C1 sky130_fd_sc_hd__o211a_1
X_10434_ VPWR VGND VPWR VGND _10433_/X _10662_/S _10667_/C1 _10434_/X sky130_fd_sc_hd__a21o_1
X_10365_ VGND VPWR VPWR VGND _10365_/X hold827/A _10604_/S hold818/A sky130_fd_sc_hd__mux2_1
X_12104_ VGND VPWR VPWR VGND _12104_/X hold800/A _12117_/B hold440/A sky130_fd_sc_hd__mux2_1
X_10296_ VGND VPWR VGND VPWR _10296_/X _15004_/Q _10633_/A2 _10295_/X _10288_/S sky130_fd_sc_hd__o211a_1
X_12035_ VGND VPWR VPWR VGND _12035_/X _14874_/Q _12112_/S hold361/A sky130_fd_sc_hd__mux2_1
XFILLER_26_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_24_1261 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_1366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_1379 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12868_ VGND VPWR VPWR VGND _15592_/D _12868_/A1 _12870_/S _15592_/Q sky130_fd_sc_hd__mux2_1
X_11819_ VGND VPWR VGND VPWR _11819_/X _11816_/X _11818_/X _12748_/A1 _12748_/C1 sky130_fd_sc_hd__a211o_1
X_14607_ hold746/A _14607_/CLK _14607_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15587_ _15587_/Q clkload44/A _15587_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12799_ VPWR VGND VGND VPWR _12799_/X _12822_/A _12799_/B sky130_fd_sc_hd__or2_1
X_14538_ _14538_/Q _14538_/CLK _14538_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14469_ hold658/A _14469_/CLK _14469_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13112__229 VPWR VGND VPWR VGND _14355_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_12982__99 VPWR VGND VPWR VGND _14225_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_08961_ VGND VPWR VGND VPWR _15117_/D hold985/X _08985_/A2 _08960_/X _08955_/A sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_65_Right_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13463__580 VPWR VGND VPWR VGND _14738_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_07912_ VGND VPWR VGND VPWR _07912_/X _15140_/Q _15351_/Q clone13/A clone18/A sky130_fd_sc_hd__a22o_4
X_08892_ VPWR VGND VGND VPWR _08892_/X _15146_/Q _08918_/B sky130_fd_sc_hd__or2_1
X_07843_ VPWR VGND VGND VPWR _15564_/Q _07885_/A _07906_/A sky130_fd_sc_hd__nand2_1
X_13006__123 VPWR VGND VPWR VGND _14249_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
XFILLER_77_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07774_ VGND VPWR VGND VPWR _08218_/B _07773_/B _08247_/A _07773_/A sky130_fd_sc_hd__a21bo_1
X_09513_ VGND VPWR VPWR VGND _14546_/D _09860_/A0 _09513_/S hold665/X sky130_fd_sc_hd__mux2_1
XFILLER_77_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13810__927 VPWR VGND VPWR VGND _15182_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_09444_ VGND VPWR VPWR VGND _14608_/D _09862_/A0 _09449_/S hold784/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_74_Right_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09375_ VGND VPWR VPWR VGND _14671_/D hold638/X _09376_/S _09829_/A1 sky130_fd_sc_hd__mux2_1
X_08326_ VGND VPWR VPWR VGND _15493_/D fanout17/X _08338_/S hold844/X sky130_fd_sc_hd__mux2_1
X_08257_ VGND VPWR VPWR VGND _10061_/A _08257_/X _08257_/B sky130_fd_sc_hd__xor2_1
XFILLER_14_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08188_ VPWR VGND VGND VPWR _07993_/A _08186_/Y _08220_/A _08187_/Y _08188_/X sky130_fd_sc_hd__o22a_1
X_07208_ VGND VPWR VPWR VGND _07230_/S _15596_/Q _14385_/Q _07372_/C sky130_fd_sc_hd__mux2_2
Xclkbuf_3_5_0_clk clkload3/A clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07139_ VGND VPWR VGND VPWR _15574_/Q _07141_/A _07827_/D sky130_fd_sc_hd__or2_4
XFILLER_3_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13704__821 VPWR VGND VPWR VGND _15044_/CLK clkload16/A sky130_fd_sc_hd__inv_2
X_10150_ VGND VPWR VPWR VGND _10150_/X hold498/A _10604_/S hold727/A sky130_fd_sc_hd__mux2_1
X_10081_ VPWR VGND VPWR VGND _10079_/X _10060_/A _14153_/Q _10081_/Y sky130_fd_sc_hd__a21oi_1
X_14073__1190 VPWR VGND VPWR VGND _15492_/CLK clkload11/A sky130_fd_sc_hd__inv_2
XFILLER_0_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10983_ VPWR VGND VGND VPWR _10983_/X _10985_/S _10983_/B sky130_fd_sc_hd__or2_1
X_12722_ VPWR VGND VPWR VGND _12721_/X _12722_/A1 _12720_/X _12722_/Y sky130_fd_sc_hd__a21oi_1
X_15510_ hold959/A _15510_/CLK _15510_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15441_ _15441_/Q clkload47/A _15441_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_43_587 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12653_ VPWR VGND VGND VPWR _12653_/X _12655_/S _12653_/B sky130_fd_sc_hd__or2_1
X_12584_ VPWR VGND VGND VPWR _12584_/A _12584_/B _12584_/Y sky130_fd_sc_hd__nor2_1
X_15372_ hold398/A _15372_/CLK _15372_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11604_ VPWR VGND VGND VPWR _11585_/Y _11603_/X _10710_/B _15445_/Q _15445_/D _11296_/A
+ sky130_fd_sc_hd__o221a_1
X_14323_ hold884/A _14323_/CLK _14323_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11535_ VGND VPWR _11535_/X _15096_/Q _11535_/A _11535_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14254_ hold492/A _14254_/CLK _14254_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11466_ VGND VPWR VPWR VGND _11466_/X _15074_/Q _11475_/S _15072_/Q sky130_fd_sc_hd__mux2_1
X_11397_ VPWR VGND VPWR VGND _11396_/X _14852_/Q _11395_/X _14852_/D _11361_/X sky130_fd_sc_hd__a22o_1
X_14185_ hold594/A _14185_/CLK _14185_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10417_ VGND VPWR VPWR VGND _10417_/X _14484_/Q _10735_/S hold453/A sky130_fd_sc_hd__mux2_1
X_13447__564 VPWR VGND VPWR VGND _14722_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_10348_ VGND VPWR VPWR VGND _10348_/X _10345_/X _10685_/S _10344_/X sky130_fd_sc_hd__mux2_1
X_10279_ VGND VPWR VPWR VGND _10279_/X hold434/A _10602_/S hold390/A sky130_fd_sc_hd__mux2_1
X_12018_ VGND VPWR VPWR VGND _12018_/X _12015_/X _12106_/S _12014_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_1152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07490_ VPWR VGND VGND VPWR _08603_/A _08603_/B _07462_/A _08598_/A sky130_fd_sc_hd__o21a_1
X_15639_ VGND VPWR VPWR VGND _15639_/Q _15639_/D _10060_/Y sky130_fd_sc_hd__dlxtn_2
XFILLER_9_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09160_ VGND VPWR VPWR VGND _14938_/D _09228_/A0 _09160_/S hold967/X sky130_fd_sc_hd__mux2_1
X_14097__1214 VPWR VGND VPWR VGND _15516_/CLK clkload37/A sky130_fd_sc_hd__inv_2
X_08111_ VGND VPWR VGND VPWR _11302_/A _14859_/Q _08112_/A _08110_/X sky130_fd_sc_hd__a21oi_2
X_09091_ VGND VPWR VPWR VGND _15002_/D hold1111/X _09091_/S _09228_/A0 sky130_fd_sc_hd__mux2_1
X_08042_ VGND VPWR _08042_/B _12794_/B _08047_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold912 hold912/X hold912/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold901 hold901/X hold901/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 hold923/X hold923/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 hold945/X hold945/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 hold934/X hold934/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 hold989/X hold989/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ VPWR VGND VGND VPWR _15612_/Q _09993_/B _09994_/B sky130_fd_sc_hd__nor2_1
Xhold978 hold978/X hold978/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 hold956/X hold956/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 hold967/X hold967/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ VPWR VGND VPWR VGND _08972_/A _15124_/Q _08933_/A _08945_/B hold1425/X sky130_fd_sc_hd__a22o_1
XFILLER_44_1412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08875_ VGND VPWR VGND VPWR _15155_/D hold1171/X _08919_/A2 _08874_/X _11308_/C1
+ sky130_fd_sc_hd__o211a_1
X_07826_ _07826_/X _15576_/Q _07826_/A _15572_/Q _07826_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_13240__357 VPWR VGND VPWR VGND _14515_/CLK clkload19/A sky130_fd_sc_hd__inv_2
X_07757_ VGND VPWR _07777_/A _15595_/Q _15548_/Q _07757_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_53_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07688_ VPWR VGND VGND VPWR _07688_/X _07688_/A _07688_/B sky130_fd_sc_hd__or2_1
X_13093__210 VPWR VGND VPWR VGND _14336_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_13982__1099 VPWR VGND VPWR VGND _15354_/CLK clkload23/A sky130_fd_sc_hd__inv_2
X_09427_ VGND VPWR VPWR VGND _14625_/D _09446_/S clone46/A hold1248/X sky130_fd_sc_hd__mux2_4
X_09358_ VGND VPWR VPWR VGND _14688_/D hold697/X _09376_/S fanout50/X sky130_fd_sc_hd__mux2_1
X_08309_ VGND VPWR VPWR VGND _15510_/D fanout80/X _08318_/S hold959/X sky130_fd_sc_hd__mux2_1
X_11320_ VPWR VGND VGND VPWR _14826_/Q _11320_/Y _14825_/Q sky130_fd_sc_hd__nand2_1
X_09289_ VGND VPWR VPWR VGND _09307_/S fanout48/X hold1168/X _14752_/D sky130_fd_sc_hd__mux2_2
X_13134__251 VPWR VGND VPWR VGND _14377_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_11251_ VPWR VGND VGND VPWR _11251_/X _14925_/Q _11251_/B sky130_fd_sc_hd__or2_1
X_10202_ VGND VPWR VPWR VGND _10206_/B hold673/A _10567_/S hold253/A sky130_fd_sc_hd__mux2_1
X_11182_ VGND VPWR VPWR VGND _11182_/X hold657/A _11186_/S hold294/A sky130_fd_sc_hd__mux2_1
X_10133_ VGND VPWR VGND VPWR _10133_/X _10347_/A1 _10129_/X _10132_/X _10622_/C1 sky130_fd_sc_hd__o211a_1
X_14941_ hold975/A _14941_/CLK _14941_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10064_ VPWR VGND VPWR VGND _10064_/B _10064_/D _10064_/C _10064_/A _10064_/X sky130_fd_sc_hd__or4_1
X_14872_ hold781/A _14872_/CLK _14872_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_48_668 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_498 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_1325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_690 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_29_893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12998__115 VPWR VGND VPWR VGND _14241_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
XFILLER_44_863 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_1369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10966_ VGND VPWR VGND VPWR _10966_/X _15022_/Q _11252_/A2 _10965_/X _11143_/S sky130_fd_sc_hd__o211a_1
X_12705_ VGND VPWR VGND VPWR _12705_/X _15396_/Q _12705_/A2 _12748_/A1 _12704_/X sky130_fd_sc_hd__o211a_1
X_10897_ VGND VPWR VPWR VGND _10901_/B _14625_/Q _10919_/S hold450/A sky130_fd_sc_hd__mux2_1
X_15424_ hold310/A _15424_/CLK _15424_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12636_ VGND VPWR VGND VPWR _12636_/X hold930/A _12743_/A2 _12737_/B1 _12635_/X sky130_fd_sc_hd__o211a_1
XFILLER_15_1002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15355_ _15355_/Q _15355_/CLK _15355_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12567_ VGND VPWR VPWR VGND _12571_/B _14630_/Q _12578_/S _14662_/Q sky130_fd_sc_hd__mux2_1
X_14306_ hold339/A _14306_/CLK _14306_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15286_ hold950/A _15286_/CLK _15286_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11518_ VGND VPWR VPWR VGND _11518_/X _11517_/X _11537_/S _15470_/Q sky130_fd_sc_hd__mux2_1
X_12498_ VGND VPWR VGND VPWR _12498_/X _12670_/A1 _12494_/X _12497_/X _12670_/C1 sky130_fd_sc_hd__o211a_1
Xhold208 hold208/X hold208/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ hold505/A _14237_/CLK _14237_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11449_ VGND VPWR VPWR VGND _11449_/X _11448_/X _11476_/S _15447_/Q sky130_fd_sc_hd__mux2_1
Xhold219 hold219/X hold219/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13681__798 VPWR VGND VPWR VGND _15021_/CLK clkload36/A sky130_fd_sc_hd__inv_2
XFILLER_67_1445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12952__69 VPWR VGND VPWR VGND _14195_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_14168_ hold820/A _14168_/CLK _14168_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08660_ VPWR VGND VGND VPWR _08660_/X _14388_/Q _08664_/B sky130_fd_sc_hd__or2_1
XFILLER_54_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_616 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07611_ VPWR VGND VPWR VGND _15095_/Q _07881_/A2 _07611_/X _07668_/B _07154_/A _07610_/Y
+ sky130_fd_sc_hd__a221o_1
X_08591_ VPWR VGND VGND VPWR _15551_/Q _08591_/Y _08591_/B sky130_fd_sc_hd__nand2_1
X_13575__692 VPWR VGND VPWR VGND _14906_/CLK clkload10/A sky130_fd_sc_hd__inv_2
X_07542_ VPWR VGND _07542_/X _07515_/A _07513_/X _07512_/A _07523_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_50_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07473_ VGND VPWR VPWR VGND _07477_/S _12855_/A0 _15592_/Q _07482_/B sky130_fd_sc_hd__mux2_2
X_09212_ VGND VPWR VPWR VGND _14881_/D _09228_/S hold1200/X clone44/X sky130_fd_sc_hd__mux2_4
X_13118__235 VPWR VGND VPWR VGND _14361_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_09143_ VGND VPWR VPWR VGND _14955_/D fanout44/X _09160_/S hold817/X sky130_fd_sc_hd__mux2_1
X_09074_ VGND VPWR VPWR VGND _15019_/D hold1055/X _09088_/S fanout44/X sky130_fd_sc_hd__mux2_1
Xhold720 hold720/X hold720/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08025_ VGND VPWR _08025_/B _12799_/B _08025_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold742 hold742/X hold742/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 hold764/X hold764/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 hold731/X hold731/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 hold753/X hold753/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 hold786/X hold786/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 hold797/X hold797/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 hold775/X hold775/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ VPWR VGND VGND VPWR _09976_/B _12878_/C _10056_/A sky130_fd_sc_hd__nand2_4
X_08927_ VGND VPWR VGND VPWR _15129_/D input2/X _08902_/B _08926_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
X_08858_ VPWR VGND VGND VPWR _14144_/Q _08859_/C _08858_/Y sky130_fd_sc_hd__nor2_1
Xhold1420 hold1420/X _15316_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 hold1442/X _14146_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1431 hold1431/X _15588_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13816__933 VPWR VGND VPWR VGND _15188_/CLK clkload38/A sky130_fd_sc_hd__inv_2
Xhold1464 _08882_/A _15151_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07809_ VGND VPWR _07809_/B _07810_/B _07809_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold1453 hold1453/X _15278_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08789_ VGND VPWR VPWR VGND _15220_/D fanout66/X _08808_/S hold205/X sky130_fd_sc_hd__mux2_1
X_10820_ VPWR VGND VPWR VGND _10820_/X _11173_/A _10793_/X _10801_/X _10819_/X _10818_/X
+ sky130_fd_sc_hd__o32a_1
X_10751_ VGND VPWR VPWR VGND _10751_/X hold690/A _10835_/B hold182/A sky130_fd_sc_hd__mux2_1
X_10682_ VGND VPWR VGND VPWR _10682_/X _10693_/B1 _10677_/X _10681_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_12421_ VGND VPWR VPWR VGND _12421_/X hold713/A _12661_/S _15250_/Q sky130_fd_sc_hd__mux2_1
X_15140_ _15140_/Q _15140_/CLK _15140_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12352_ VGND VPWR VGND VPWR _12352_/X _12351_/X _12350_/X _12367_/S _12863_/A1 sky130_fd_sc_hd__a211o_1
X_11303_ VPWR VGND VGND VPWR _11303_/A _11303_/Y _11303_/B sky130_fd_sc_hd__nand2_1
X_12283_ VPWR VGND VGND VPWR _12283_/X _12698_/S _12283_/B sky130_fd_sc_hd__or2_1
X_15071_ _15071_/Q clkload15/A _15071_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11234_ VPWR VGND VGND VPWR _11234_/X _11244_/S _11234_/B sky130_fd_sc_hd__or2_1
XFILLER_5_778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11165_ VGND VPWR VPWR VGND _11165_/X hold535/A _11165_/S hold262/A sky130_fd_sc_hd__mux2_1
X_11096_ VGND VPWR VGND VPWR _11096_/X _11093_/X _11095_/X _11215_/C1 _11096_/C1 sky130_fd_sc_hd__a211o_1
X_14096__1213 VPWR VGND VPWR VGND _15515_/CLK clkload22/A sky130_fd_sc_hd__inv_2
XFILLER_0_461 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10116_ VGND VPWR VGND VPWR _10116_/X _10113_/X _10115_/X _10614_/A1 _10608_/A1 sky130_fd_sc_hd__a211o_1
XFILLER_48_421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10047_ VPWR VGND VGND VPWR _10049_/B _10047_/B _15635_/D sky130_fd_sc_hd__nor2_1
X_14924_ hold329/A _14924_/CLK _14924_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_76_796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_36_616 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13559__676 VPWR VGND VPWR VGND _14890_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
X_14855_ _14855_/Q clkload26/A _14855_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14786_ hold493/A _14786_/CLK _14786_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11998_ VGND VPWR VPWR VGND _11998_/X hold994/A _11998_/S hold650/A sky130_fd_sc_hd__mux2_1
XFILLER_44_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_671 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10949_ VPWR VGND VPWR VGND _10948_/X _11181_/A1 _10947_/X _10949_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_1168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14052__1169 VPWR VGND VPWR VGND _15424_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_15407_ hold612/A _15407_/CLK _15407_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12619_ VPWR VGND VPWR VGND _12618_/X _12740_/A1 _12617_/X _12619_/Y sky130_fd_sc_hd__a21oi_1
X_15338_ _15338_/Q _15338_/CLK _15338_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15269_ _15269_/Q _15269_/CLK _15269_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14191__909 _14191_/D _14191__909/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xfanout529 VGND VPWR _12594_/B _12589_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13981__1098 VPWR VGND VPWR VGND _15353_/CLK clkload23/A sky130_fd_sc_hd__inv_2
XFILLER_59_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13503__620 VPWR VGND VPWR VGND _14778_/CLK _12954__71/A sky130_fd_sc_hd__inv_2
X_09830_ VGND VPWR VPWR VGND _14222_/D _09864_/A0 _09830_/S hold253/X sky130_fd_sc_hd__mux2_1
Xfanout518 VGND VPWR _12446_/B _12635_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout507 VGND VPWR _12477_/B _12479_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_80_1453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09761_ VGND VPWR VPWR VGND _14285_/D _09865_/A0 _09763_/S hold278/X sky130_fd_sc_hd__mux2_1
XFILLER_67_741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_41_1426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08712_ VGND VPWR VGND VPWR _08712_/X _08714_/A2 _08726_/C1 hold982/X _08711_/X sky130_fd_sc_hd__a211o_1
Xrebuffer12 VPWR VGND VPWR VGND _09486_/A _15578_/Q sky130_fd_sc_hd__dlygate4sd1_1
X_09692_ VGND VPWR VPWR VGND _14348_/D hold871/X _09693_/S _09692_/A0 sky130_fd_sc_hd__mux2_1
Xrebuffer23 VPWR VGND VPWR VGND rebuffer23/X rebuffer24/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer34 VPWR VGND VPWR VGND rebuffer34/X rebuffer35/X sky130_fd_sc_hd__dlygate4sd1_1
X_08643_ VGND VPWR VGND VPWR _15297_/D hold1035/X _08704_/A2 _08642_/X _11937_/C1
+ sky130_fd_sc_hd__o211a_1
X_08574_ VPWR VGND VPWR VGND _08580_/B _08580_/A _07450_/A _08575_/B sky130_fd_sc_hd__a21oi_1
XFILLER_54_468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07525_ VPWR VGND _07526_/B _07519_/Y _07518_/X _07429_/A _08604_/B2 VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_35_1219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clk clkload17/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_07456_ VPWR VGND VPWR VGND _07455_/X _07447_/A _07454_/X _07456_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13352__469 VPWR VGND VPWR VGND _14627_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_07387_ VGND VPWR VGND VPWR _07387_/X _08007_/A _07982_/B _07389_/B sky130_fd_sc_hd__a21bo_1
X_09126_ VGND VPWR VPWR VGND _14969_/D hold777/X _09126_/S _09691_/A0 sky130_fd_sc_hd__mux2_1
X_09057_ VGND VPWR VPWR VGND _15033_/D hold653/X _09059_/S _09691_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_11_1241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08008_ VPWR VGND _08008_/X _10065_/B _08182_/S VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_2_704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold572 hold572/X hold572/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 hold561/X hold561/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 hold550/X hold550/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 hold594/X hold594/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13246__363 VPWR VGND VPWR VGND _14521_/CLK clkload10/A sky130_fd_sc_hd__inv_2
Xhold583 hold583/X hold583/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09959_ _14803_/D _15259_/Q _15063_/Q _14804_/Q _08591_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_79_1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold1261 hold1261/X _15156_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1250 _15154_/D _08877_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1294 hold1294/X _15149_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1283 _15363_/D _08427_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 hold1272/X _15600_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ VGND VPWR VPWR VGND _11921_/X hold525/A _12149_/S hold644/A sky130_fd_sc_hd__mux2_1
XFILLER_45_457 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11852_ VGND VPWR VGND VPWR _11852_/X _12008_/C1 _11847_/X _11851_/X _12111_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_2_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14640_ hold449/A _14640_/CLK _14640_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10803_ VGND VPWR VPWR VGND _10803_/X hold852/A _11216_/S hold762/A sky130_fd_sc_hd__mux2_1
X_14571_ hold199/A _14571_/CLK _14571_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clkload34/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_11783_ VGND VPWR VPWR VGND _11783_/X hold523/A _12205_/S hold555/A sky130_fd_sc_hd__mux2_1
XFILLER_40_162 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10734_ VGND VPWR VGND VPWR _10734_/X hold792/A _10744_/A2 _10733_/X _10745_/A1 sky130_fd_sc_hd__o211a_1
X_10665_ VPWR VGND VGND VPWR _10665_/X hold457/A _10670_/S sky130_fd_sc_hd__or2_1
X_12404_ VGND VPWR VGND VPWR _12404_/X hold831/A _12488_/A2 _12720_/A1 _12403_/X sky130_fd_sc_hd__o211a_1
X_15123_ _15123_/Q _15123_/CLK _15123_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12335_ VPWR VGND VGND VPWR _12335_/X hold228/A _12339_/B sky130_fd_sc_hd__or2_1
X_10596_ VGND VPWR VGND VPWR _10596_/X _15012_/Q _10744_/A2 _10595_/X _10588_/S sky130_fd_sc_hd__o211a_1
X_12266_ VGND VPWR VPWR VGND _12266_/X _12265_/X _12583_/S _12257_/X sky130_fd_sc_hd__mux2_1
X_15054_ hold346/A _15054_/CLK _15054_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12922__39 VPWR VGND VPWR VGND _14165_/CLK clkload22/A sky130_fd_sc_hd__inv_2
X_11217_ VGND VPWR VGND VPWR _11217_/X _11216_/X _11215_/X _11213_/S _11217_/C1 sky130_fd_sc_hd__a211o_1
X_12197_ VGND VPWR VPWR VGND _12201_/B hold618/A _12228_/B hold319/A sky130_fd_sc_hd__mux2_1
X_11148_ VGND VPWR VGND VPWR _11148_/X _11145_/X _11147_/X _11189_/A1 _11254_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_49_763 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11079_ VPWR VGND _11079_/X _11078_/X _11074_/X _11246_/S _11070_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14907_ hold298/A _14907_/CLK _14907_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14838_ _14838_/Q clkload28/A _14838_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_52_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07310_ VPWR VGND VPWR VGND _07298_/A _07293_/B _07291_/X _07310_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_43_clk clkload33/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_14769_ hold427/A _14769_/CLK _14769_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08290_ VGND VPWR _08290_/B _10061_/D _08290_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07241_ VPWR VGND _07241_/X _07376_/B _15454_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_13189__306 VPWR VGND VPWR VGND _14464_/CLK clkload48/A sky130_fd_sc_hd__inv_2
X_07172_ VPWR VGND _07314_/A _07173_/B _15470_/Q VPWR VGND sky130_fd_sc_hd__and2_1
Xfanout304 VGND VPWR fanout314/X _10479_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout348 VPWR VGND _10795_/S fanout349/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout326 VGND VPWR _07893_/X _11241_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09813_ VGND VPWR VPWR VGND _14239_/D fanout46/X _09827_/S hold244/X sky130_fd_sc_hd__mux2_1
XFILLER_59_505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout337 VPWR VGND _10964_/S fanout349/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout315 VGND VPWR _10972_/S _10567_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_80_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout359 VGND VPWR _08195_/C _10703_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1370 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09744_ VGND VPWR VPWR VGND _14302_/D _09760_/S fanout42/X hold1157/X sky130_fd_sc_hd__mux2_4
X_09675_ VGND VPWR VPWR VGND _14365_/D hold869/X _09675_/S fanout38/X sky130_fd_sc_hd__mux2_1
XFILLER_41_1289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08626_ VPWR VGND VGND VPWR _08626_/A _10060_/C _08626_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_928 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_42_416 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08557_ VGND VPWR VGND VPWR _08557_/X _08605_/A _08627_/C1 hold905/X _08556_/Y sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_34_clk clkload52/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_70_747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08488_ VPWR VGND VGND VPWR _08488_/X _15332_/Q _08488_/B sky130_fd_sc_hd__or2_1
X_07508_ _07530_/C _07545_/A _07509_/C _07531_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_07439_ VPWR VGND VGND VPWR _15459_/Q _07507_/B _07440_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_471 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14095__1212 VPWR VGND VPWR VGND _15514_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_10_335 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10450_ VPWR VGND VPWR VGND _10450_/X _10729_/A _10423_/X _10431_/X _10449_/X _10448_/X
+ sky130_fd_sc_hd__o32a_1
X_09109_ VGND VPWR VPWR VGND _14986_/D hold891/X _09122_/S fanout41/X sky130_fd_sc_hd__mux2_1
X_10381_ VGND VPWR VPWR VGND _10381_/X hold884/A _10687_/B hold161/A sky130_fd_sc_hd__mux2_1
X_12120_ VPWR VGND _12120_/X _12119_/X _12115_/X _12102_/S _12111_/X VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold380 hold380/X hold380/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12051_ VGND VPWR VPWR VGND _12051_/X hold752/A _12219_/S hold220/A sky130_fd_sc_hd__mux2_1
Xhold391 hold391/X hold391/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ VPWR VGND VGND VPWR _11002_/X hold301/A _11231_/S sky130_fd_sc_hd__or2_1
X_13480__597 VPWR VGND VPWR VGND _14755_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
XFILLER_77_346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout860 VPWR VGND _08294_/B1 _08249_/B2 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_77_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout882 VPWR VGND VGND VPWR rebuffer7/A _07703_/A sky130_fd_sc_hd__buf_8
Xfanout871 VPWR VGND _11535_/A _15600_/Q VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_24_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14051__1168 VPWR VGND VPWR VGND _15423_/CLK clkload40/A sky130_fd_sc_hd__inv_2
XFILLER_58_582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_571 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1080 hold1080/X _15311_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_34_906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold1091 hold1091/X _14942_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ VGND VPWR VPWR VGND _11904_/X hold455/A _12205_/S hold330/A sky130_fd_sc_hd__mux2_1
X_14623_ hold720/A _14623_/CLK _14623_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_73_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_61_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12884_ VPWR VGND VPWR VGND _08233_/X _07574_/A _12883_/A _15605_/D sky130_fd_sc_hd__a21oi_1
XFILLER_45_265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_clk clkload32/A clkload1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_11835_ VGND VPWR VPWR VGND _11839_/B hold485/A _12171_/S hold213/A sky130_fd_sc_hd__mux2_1
XFILLER_57_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_961 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14554_ hold745/A _14554_/CLK _14554_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11766_ VGND VPWR VGND VPWR _11766_/X _12099_/A1 _11762_/X _11765_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
X_13374__491 VPWR VGND VPWR VGND _14649_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_13980__1097 VPWR VGND VPWR VGND _15352_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_14485_ _14485_/Q _14485_/CLK _14485_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10717_ VGND VPWR VGND VPWR _10717_/X _10745_/A1 _10713_/X _10716_/X _10717_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_70_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11697_ VGND VPWR VPWR VGND _11697_/X hold833/A _12052_/S hold672/A sky130_fd_sc_hd__mux2_1
Xrebuffer3 VPWR VGND VPWR VGND _07476_/B _07479_/A sky130_fd_sc_hd__dlymetal6s4s_1
X_10648_ VGND VPWR VPWR VGND _10648_/X _14202_/Q _10670_/S hold328/A sky130_fd_sc_hd__mux2_1
X_10579_ VPWR VGND VPWR VGND _10578_/X _10745_/C1 _10577_/X _10579_/Y sky130_fd_sc_hd__a21oi_1
X_12318_ VGND VPWR VPWR VGND _12318_/X _14207_/Q _12318_/S hold274/A sky130_fd_sc_hd__mux2_1
X_15106_ _15106_/Q _15106_/CLK _15106_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13721__838 VPWR VGND VPWR VGND _15061_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_12249_ VGND VPWR VGND VPWR _12249_/X _12702_/C1 _12244_/X _12248_/X _12583_/S sky130_fd_sc_hd__o211a_1
X_15037_ hold495/A _15037_/CLK _15037_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_69_836 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07790_ VPWR VGND VGND VPWR _07795_/C _07998_/C _07790_/B sky130_fd_sc_hd__nand2_1
X_09460_ VGND VPWR VPWR VGND _14596_/D fanout66/X _09467_/S hold467/X sky130_fd_sc_hd__mux2_1
X_13615__732 VPWR VGND VPWR VGND _14955_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_08411_ VGND VPWR VPWR VGND _15366_/D fanout96/X _08411_/S hold931/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_clk clkload24/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_52_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09391_ VGND VPWR VPWR VGND _14658_/D hold559/X _09408_/S clone55/X sky130_fd_sc_hd__mux2_1
X_08342_ VPWR VGND VPWR VGND _08342_/X _09729_/A _09198_/C sky130_fd_sc_hd__or2_2
X_08273_ VPWR VGND VGND VPWR _08273_/A _08273_/Y _08273_/B sky130_fd_sc_hd__nand2_1
X_14197__915 _14197_/D _14197__915/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_07224_ VPWR VGND VGND VPWR _12878_/B _07827_/C _10059_/A _07827_/A _07224_/X _07113_/Y
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_677 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07155_ VPWR VGND VGND VPWR _14408_/Q _07301_/A2 _07301_/B1 _07157_/B sky130_fd_sc_hd__o21a_1
XFILLER_3_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07086_ VPWR VGND VPWR VGND _07086_/Y _15470_/Q sky130_fd_sc_hd__inv_2
Xfanout112 VGND VPWR _08266_/X _09229_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout101 VGND VPWR _09658_/A0 _08284_/X VPWR VGND sky130_fd_sc_hd__clkbuf_1
Xfanout156 VPWR VGND _08985_/A2 _08936_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout145 VGND VPWR _08553_/A2 _08731_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout134 VPWR VGND _08722_/C1 _08726_/C1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout123 VPWR VGND _09550_/A1 _08212_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout189 VPWR VGND _12591_/S _11810_/S VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout178 VGND VPWR _07979_/X _08298_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_07988_ VPWR VGND VPWR VGND _08002_/B1 _15622_/Q _08002_/A2 _07994_/B _15586_/Q sky130_fd_sc_hd__a22o_1
Xfanout167 VGND VPWR _12106_/S _11995_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09727_ VGND VPWR VPWR VGND _14316_/D fanout99/X _09728_/S hold780/X sky130_fd_sc_hd__mux2_1
Xtt_um_femto_894 uio_oe[5] tt_um_femto_894/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_76_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_725 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13358__475 VPWR VGND VPWR VGND _14633_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_09658_ VGND VPWR VPWR VGND _14412_/D hold983/X _09659_/S _09658_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_76_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08609_ VGND VPWR VPWR VGND _08609_/A _08609_/X _08609_/B sky130_fd_sc_hd__xor2_1
X_09589_ VGND VPWR VPWR VGND _14476_/D hold1019/X _09590_/S fanout99/X sky130_fd_sc_hd__mux2_1
XFILLER_54_1414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11620_ VPWR VGND VPWR VGND _11619_/X _12008_/C1 _11618_/X _11620_/Y sky130_fd_sc_hd__a21oi_1
X_11551_ VPWR VGND VGND VPWR _11551_/A _11551_/Y _11551_/B sky130_fd_sc_hd__nand2_1
X_10502_ VPWR VGND VGND VPWR _10502_/X _10510_/S _10502_/B sky130_fd_sc_hd__or2_1
X_14270_ hold790/A _14270_/CLK _14270_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11482_ VGND VPWR VPWR VGND _11482_/X _11481_/X _11491_/S _15458_/Q sky130_fd_sc_hd__mux2_1
X_10433_ VGND VPWR VPWR VGND _10433_/X hold981/A _10553_/S hold674/A sky130_fd_sc_hd__mux2_1
X_10364_ VGND VPWR VGND VPWR _10364_/X _14942_/Q _10629_/A2 _10363_/X _10614_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_6_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_48_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_12103_ VPWR VGND VGND VPWR _12103_/A _12103_/B _12103_/Y sky130_fd_sc_hd__nor2_1
X_10295_ VPWR VGND VGND VPWR _10295_/X hold433/A _10627_/S sky130_fd_sc_hd__or2_1
X_12034_ VGND VPWR VGND VPWR _12034_/X hold637/A _12118_/A2 _12119_/A1 _12033_/X sky130_fd_sc_hd__o211a_1
Xfanout690 VPWR VGND _08332_/S _08335_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_12867_ VGND VPWR VPWR VGND _15591_/D _10333_/A _14802_/D _15591_/Q sky130_fd_sc_hd__mux2_1
X_11818_ VGND VPWR VGND VPWR _11818_/X hold782/A _12746_/A2 _12367_/S _11817_/X sky130_fd_sc_hd__o211a_1
X_15586_ _15586_/Q clkload44/A _15586_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14606_ hold368/A _14606_/CLK _14606_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12798_ VPWR VGND VGND VPWR _12822_/A _12798_/Y _12798_/B sky130_fd_sc_hd__nand2_1
X_14537_ hold210/A _14537_/CLK _14537_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11749_ VGND VPWR VGND VPWR _11749_/X _11748_/X _11747_/X _12720_/A1 _12720_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_31_1233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14468_ hold587/A _14468_/CLK _14468_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14399_ _14399_/Q clkload54/A _14399_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13151__268 VPWR VGND VPWR VGND _14426_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
X_08960_ VPWR VGND VGND VPWR _08960_/X _08969_/A _08960_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_5_clk clkload9/A clkbuf_3_0_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_08891_ VGND VPWR VGND VPWR _15147_/D hold1293/X _08893_/A2 _08890_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_07911_ VGND VPWR VPWR VGND _15533_/D fanout45/X _07954_/S hold305/X sky130_fd_sc_hd__mux2_1
X_07842_ VPWR VGND _07906_/A _07931_/A _15563_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_29_519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13045__162 VPWR VGND VPWR VGND _14288_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_14094__1211 VPWR VGND VPWR VGND _15513_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_07773_ VPWR VGND VGND VPWR _07773_/A _08247_/B _07773_/B sky130_fd_sc_hd__nand2_1
X_09512_ VGND VPWR VPWR VGND _14547_/D _09859_/A0 _09520_/S hold522/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09443_ VGND VPWR VPWR VGND _14609_/D _09827_/A1 _09443_/S hold374/X sky130_fd_sc_hd__mux2_1
XFILLER_52_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_75_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09374_ VGND VPWR VPWR VGND _14672_/D hold671/X _09379_/S _09688_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_80_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_791 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08325_ VGND VPWR VPWR VGND _15494_/D fanout21/X _08330_/S hold1028/X sky130_fd_sc_hd__mux2_1
XFILLER_32_1008 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08256_ VPWR VGND _08256_/X _08256_/B _08273_/A VPWR VGND sky130_fd_sc_hd__xor2_2
X_14050__1167 VPWR VGND VPWR VGND _15422_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_12958__75 VPWR VGND VPWR VGND _14201_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_08187_ VGND VPWR _08187_/B _08187_/Y _08187_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07207_ VGND VPWR VGND VPWR _08162_/A _07371_/B _07371_/A sky130_fd_sc_hd__xnor2_4
XFILLER_14_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13743__860 VPWR VGND VPWR VGND _15115_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_07138_ VPWR VGND VGND VPWR _15574_/Q _07826_/D _07765_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_58_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10080_ VGND VPWR VPWR VGND _10080_/X _12790_/A _08276_/Y _08273_/Y _12829_/S sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_1148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10982_ VGND VPWR VPWR VGND _10982_/X hold597/A _10994_/S hold413/A sky130_fd_sc_hd__mux2_1
XFILLER_21_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12721_ VGND VPWR VPWR VGND _12721_/X _12718_/X _12721_/S _12717_/X sky130_fd_sc_hd__mux2_1
X_15440_ _15440_/Q clkload47/A _15440_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12652_ VGND VPWR VPWR VGND _12652_/X hold656/A _12652_/S hold299/A sky130_fd_sc_hd__mux2_1
XFILLER_43_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11603_ VPWR VGND VPWR VGND _11602_/X _12103_/A _12121_/B1 _11603_/X sky130_fd_sc_hd__a21o_1
X_12583_ VGND VPWR VPWR VGND _12584_/B _12582_/Y _12583_/S _12574_/Y sky130_fd_sc_hd__mux2_1
X_15371_ hold473/A _15371_/CLK _15371_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14322_ hold761/A _14322_/CLK _14322_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11534_ VGND VPWR VPWR VGND _15095_/D _11533_/X _11538_/S _15095_/Q sky130_fd_sc_hd__mux2_1
XFILLER_7_412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_14253_ _14253_/Q _14253_/CLK _14253_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11465_ VGND VPWR VPWR VGND _15072_/D _11464_/X _11480_/S _15072_/Q sky130_fd_sc_hd__mux2_1
XFILLER_7_434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10416_ VGND VPWR VPWR VGND _10416_/X hold677/A _10720_/S hold481/A sky130_fd_sc_hd__mux2_1
X_11396_ VPWR VGND _11396_/X _11418_/S _11398_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_14184_ _14184_/Q _14184_/CLK _14184_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10347_ VGND VPWR VGND VPWR _10347_/X _10347_/A1 _10343_/X _10346_/X _10614_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_79_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13792__909 VPWR VGND VPWR VGND _15164_/CLK clkload7/A sky130_fd_sc_hd__inv_2
XFILLER_26_1302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10278_ VGND VPWR VPWR VGND _10278_/X _14192_/Q _10609_/S hold404/A sky130_fd_sc_hd__mux2_1
X_13029__146 VPWR VGND VPWR VGND _14272_/CLK clkload46/A sky130_fd_sc_hd__inv_2
XFILLER_39_817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12017_ VGND VPWR VGND VPWR _12017_/X _12119_/A1 _12013_/X _12016_/X _12017_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_26_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13686__803 VPWR VGND VPWR VGND _15026_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_15638_ VGND VPWR VPWR VGND _15638_/Q _15638_/D _10060_/Y sky130_fd_sc_hd__dlxtn_2
X_15569_ _15569_/Q clkload16/A _15569_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08110_ VPWR VGND VPWR VGND _08252_/A2 _15341_/Q _08253_/A2 _08110_/X _15146_/Q sky130_fd_sc_hd__a22o_1
X_09090_ VGND VPWR VPWR VGND _15003_/D hold1094/X _09090_/S _09689_/A0 sky130_fd_sc_hd__mux2_1
X_13727__844 VPWR VGND VPWR VGND _15099_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_08041_ VPWR VGND VGND VPWR _08041_/A _08041_/B _08042_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_1074 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold902 hold902/X hold902/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 hold913/X hold913/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 hold924/X hold924/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 hold946/X hold946/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 hold935/X hold935/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 hold957/X hold957/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold979 hold979/X hold979/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ VPWR VGND _09996_/C _09993_/B _15612_/Q VPWR VGND sky130_fd_sc_hd__and2_1
Xhold968 hold968/X hold968/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ VPWR VGND _15126_/D _08943_/B _08943_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_44_1424 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08874_ VPWR VGND VGND VPWR _08874_/X _08874_/A _08918_/B sky130_fd_sc_hd__or2_1
X_07825_ _07849_/B _07822_/X _07823_/X _07824_/X _08249_/B2 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_07756_ _08187_/A _07754_/X _07756_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_77_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07687_ VPWR VGND VPWR VGND _15631_/Q _07952_/A2 _07688_/B _07908_/B1 _15595_/Q _07686_/X
+ sky130_fd_sc_hd__a221o_1
X_09426_ VGND VPWR VPWR VGND _14626_/D fanout56/X _09443_/S hold567/X sky130_fd_sc_hd__mux2_1
XFILLER_53_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09357_ VGND VPWR VPWR VGND _14689_/D _09357_/S hold1184/X clone46/X sky130_fd_sc_hd__mux2_4
X_08308_ VGND VPWR VPWR VGND _15511_/D fanout83/X _08318_/S hold814/X sky130_fd_sc_hd__mux2_1
X_09288_ VGND VPWR VPWR VGND _14753_/D _09307_/S clone46/X hold1158/X sky130_fd_sc_hd__mux2_4
X_13173__290 VPWR VGND VPWR VGND _14448_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_15264__939 _15264_/D _15264__939/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08239_ VGND VPWR _10062_/A _08240_/B _08239_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_69_23 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_1335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11250_ VGND VPWR VPWR VGND _11250_/X _11249_/X _11250_/S _11248_/X sky130_fd_sc_hd__mux2_1
X_10201_ VPWR VGND VPWR VGND _10200_/X _11237_/A1 _10199_/X _10201_/Y sky130_fd_sc_hd__a21oi_1
X_11181_ VGND VPWR VGND VPWR _11181_/X _11181_/A1 _11176_/X _11180_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
X_10132_ VPWR VGND VGND VPWR _10132_/X _10615_/S _10132_/B sky130_fd_sc_hd__or2_1
X_13520__637 VPWR VGND VPWR VGND _14795_/CLK clkload53/A sky130_fd_sc_hd__inv_2
XFILLER_47_1092 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10063_ VPWR VGND VPWR VGND _10063_/B _10063_/D _10063_/C _10063_/A _10064_/D sky130_fd_sc_hd__or4_1
X_14940_ hold856/A _14940_/CLK _14940_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14871_ _14871_/Q _14871_/CLK _14871_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_1337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12704_ VPWR VGND VGND VPWR _12704_/X hold325/A _12708_/S sky130_fd_sc_hd__or2_1
X_10965_ VPWR VGND VGND VPWR _10965_/X hold471/A _11142_/S sky130_fd_sc_hd__or2_1
X_10896_ VGND VPWR VGND VPWR _14400_/D _12491_/B1 _10894_/X _10895_/X _07544_/B sky130_fd_sc_hd__o211a_1
X_15423_ hold371/A _15423_/CLK _15423_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13414__531 VPWR VGND VPWR VGND _14689_/CLK clkload34/A sky130_fd_sc_hd__inv_2
X_12635_ VPWR VGND VGND VPWR _12635_/X hold164/A _12635_/B sky130_fd_sc_hd__or2_1
X_15354_ _15354_/Q _15354_/CLK _15354_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12566_ VPWR VGND VGND VPWR _12547_/Y _12565_/X _12751_/A2 _15471_/Q _15471_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
X_14093__1210 VPWR VGND VPWR VGND _15512_/CLK clkload54/A sky130_fd_sc_hd__inv_2
X_11517_ VGND VPWR VPWR VGND _11517_/X _15091_/Q _11529_/S _15089_/Q sky130_fd_sc_hd__mux2_1
X_14305_ _14305_/Q _14305_/CLK _14305_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15285_ _15285_/Q _15285_/CLK _15285_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12497_ VPWR VGND VGND VPWR _12497_/X _12665_/S _12497_/B sky130_fd_sc_hd__or2_1
Xhold209 hold209/X hold209/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ VGND VPWR VPWR VGND _11448_/X _15068_/Q _11475_/S _15066_/Q sky130_fd_sc_hd__mux2_1
X_14236_ hold334/A _14236_/CLK _14236_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11379_ VGND VPWR VPWR VGND _14846_/D _11378_/X _11382_/S hold1296/X sky130_fd_sc_hd__mux2_1
X_14167_ hold848/A _14167_/CLK _14167_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_79_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1007 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08590_ VGND VPWR VGND VPWR _15309_/D hold989/X _08628_/A2 _08589_/X _09000_/C1 sky130_fd_sc_hd__o211a_1
X_07610_ VPWR VGND VGND VPWR _07610_/A _07972_/B _07610_/Y sky130_fd_sc_hd__nor2_1
X_07541_ VPWR VGND VPWR VGND _07513_/X _07512_/A _07515_/A _07541_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_3_4_0_clk clkload2/A clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_19_393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07472_ VPWR VGND VPWR VGND _07577_/B _07486_/B sky130_fd_sc_hd__inv_2
X_13157__274 VPWR VGND VPWR VGND _14432_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_09211_ VGND VPWR VPWR VGND _14882_/D hold846/X _09228_/S fanout44/X sky130_fd_sc_hd__mux2_1
X_09142_ VGND VPWR VPWR VGND _14956_/D _09160_/S fanout50/X hold1247/X sky130_fd_sc_hd__mux2_4
X_09073_ VGND VPWR VPWR VGND _15020_/D hold1053/X _09090_/S clone100/X sky130_fd_sc_hd__mux2_1
X_12928__45 VPWR VGND VPWR VGND _14171_/CLK clkload21/A sky130_fd_sc_hd__inv_2
XFILLER_11_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold710 hold710/X hold710/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08024_ VPWR VGND VGND VPWR _08220_/A _08020_/Y _07993_/A _08023_/X _08024_/X sky130_fd_sc_hd__o22a_1
Xhold721 hold721/X hold721/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 hold743/X hold743/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 hold754/X hold754/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 hold732/X hold732/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 hold787/X hold787/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 hold776/X hold776/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 hold765/X hold765/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ VPWR VGND VGND VPWR _09975_/A _11340_/A _09975_/Y sky130_fd_sc_hd__nor2_1
Xhold798 hold798/X hold798/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ VPWR VGND VGND VPWR _08926_/X _15129_/Q _08926_/B sky130_fd_sc_hd__or2_1
Xhold1410 hold1410/X _15030_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08857_ VPWR VGND VPWR VGND _08857_/Y _08859_/C sky130_fd_sc_hd__inv_2
Xhold1421 hold1421/X _15328_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 hold1432/X _15127_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 hold1443/X hold928/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13855__972 VPWR VGND VPWR VGND _15227_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_24_Left_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1454 _08466_/A _15343_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07808_ VGND VPWR _07808_/B _07809_/B _15566_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold1465 hold1465/X hold953/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08788_ VGND VPWR VPWR VGND _15221_/D fanout70/X _08808_/S hold285/X sky130_fd_sc_hd__mux2_1
X_07739_ VPWR VGND VGND VPWR _08056_/B _15555_/Q _07739_/B sky130_fd_sc_hd__or2_1
X_10750_ VGND VPWR VPWR VGND _10750_/X _14493_/Q _10835_/B hold855/A sky130_fd_sc_hd__mux2_1
X_10681_ VGND VPWR VGND VPWR _10681_/X _10680_/X _10679_/X _10685_/S _10697_/B1 sky130_fd_sc_hd__a211o_1
XFILLER_41_845 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09409_ VGND VPWR VPWR VGND _14640_/D hold449/X _09414_/S _09723_/A1 sky130_fd_sc_hd__mux2_1
XFILLER_71_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_51_1203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12420_ VGND VPWR VPWR VGND _12420_/X hold787/A _12661_/S hold825/A sky130_fd_sc_hd__mux2_1
X_12351_ VGND VPWR VPWR VGND _12351_/X _14560_/Q _12370_/S hold254/A sky130_fd_sc_hd__mux2_1
X_11302_ VPWR VGND VGND VPWR _11302_/A _11303_/B _11302_/B sky130_fd_sc_hd__nand2_1
X_12282_ VGND VPWR VPWR VGND _12282_/X hold378/A _12282_/S hold620/A sky130_fd_sc_hd__mux2_1
X_15070_ _15070_/Q clkload15/A _15070_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11233_ VGND VPWR VPWR VGND _11233_/X _14570_/Q _11240_/S _14602_/Q sky130_fd_sc_hd__mux2_1
X_11164_ VGND VPWR VPWR VGND _11168_/B hold732/A _11167_/S hold276/A sky130_fd_sc_hd__mux2_1
X_11095_ VGND VPWR VGND VPWR _11095_/X _14278_/Q _11262_/A2 _11094_/X _11092_/S sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_42_Left_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10115_ VGND VPWR VGND VPWR _10115_/X _14999_/Q _10629_/A2 _10114_/X _10144_/S sky130_fd_sc_hd__o211a_1
X_10046_ VPWR VGND VPWR VGND _10045_/C hold1457/X hold1281/X _10047_/B sky130_fd_sc_hd__a21oi_1
X_14923_ hold424/A _14923_/CLK _14923_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14854_ _14854_/Q clkload26/A _14854_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14785_ hold749/A _14785_/CLK _14785_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11997_ VGND VPWR VGND VPWR _11997_/X _14946_/Q _12188_/A2 _12008_/A1 _11996_/X sky130_fd_sc_hd__o211a_1
X_10948_ VGND VPWR VPWR VGND _10948_/X _10945_/X _11170_/S _10944_/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_51_Left_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10879_ VPWR VGND VPWR VGND _10876_/X _10890_/A _10878_/X _10879_/X sky130_fd_sc_hd__a21o_1
X_15406_ hold725/A _15406_/CLK _15406_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1423 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12618_ VGND VPWR VPWR VGND _12618_/X _12615_/X _12624_/S _12614_/X sky130_fd_sc_hd__mux2_1
X_15337_ _15337_/Q _15337_/CLK _15337_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12549_ VGND VPWR VGND VPWR _12549_/X hold935/A _12669_/A2 _12665_/S _12548_/X sky130_fd_sc_hd__o211a_1
XFILLER_8_551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XANTENNA_1 _07561_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_15268_ _15268_/Q _15268_/CLK _15268_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13798__915 VPWR VGND VPWR VGND _15170_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_14219_ hold320/A _14219_/CLK _14219_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15199_ hold264/A _15199_/CLK _15199_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_60_Left_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout519 VGND VPWR _12446_/B _12736_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout508 VPWR VGND _12477_/B _12716_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_13839__956 VPWR VGND VPWR VGND _15211_/CLK clkload21/A sky130_fd_sc_hd__inv_2
X_09760_ VGND VPWR VPWR VGND _14286_/D _09864_/A0 _09760_/S hold259/X sky130_fd_sc_hd__mux2_1
X_09691_ VGND VPWR VPWR VGND _14349_/D hold1023/X _09693_/S _09691_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_41_1438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_444 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08711_ VGND VPWR VGND VPWR _08711_/X _14388_/Q _08664_/B _08711_/B1 _08659_/Y sky130_fd_sc_hd__o211a_1
X_08642_ VPWR VGND VPWR VGND hold907/A _08667_/A2 _08642_/X _08662_/B1 _08641_/X _08700_/B1
+ sky130_fd_sc_hd__a221o_1
Xrebuffer35 VPWR VGND VPWR VGND rebuffer35/X rebuffer36/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer24 VPWR VGND VPWR VGND rebuffer24/X rebuffer25/X sky130_fd_sc_hd__dlygate4sd1_1
X_08573_ VPWR VGND VGND VPWR _07494_/X _15599_/Q _15454_/Q _07453_/X _08580_/B sky130_fd_sc_hd__o22a_1
X_07524_ VPWR VGND VGND VPWR _08943_/A _07524_/Y _07534_/B sky130_fd_sc_hd__nand2_1
X_07455_ VPWR VGND VPWR VGND _07714_/A _15456_/Q _07450_/A _07455_/X sky130_fd_sc_hd__a21o_1
XFILLER_62_491 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07386_ _07389_/B _07925_/A _07971_/A _07981_/A _07945_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_09125_ VGND VPWR VPWR VGND _14970_/D hold406/X _09125_/S _09228_/A0 sky130_fd_sc_hd__mux2_1
X_09056_ VGND VPWR VPWR VGND _15034_/D hold614/X _09056_/S _09228_/A0 sky130_fd_sc_hd__mux2_1
X_08007_ VPWR VGND VGND VPWR _08007_/A _10065_/B _08007_/B sky130_fd_sc_hd__nand2_1
X_13949__1066 VPWR VGND VPWR VGND _15321_/CLK clkload26/A sky130_fd_sc_hd__inv_2
Xhold551 hold551/X hold551/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 hold562/X hold562/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_716 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xhold540 hold540/X hold540/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold573/X hold573/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 hold584/X hold584/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold595/X hold595/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09958_ VPWR VGND VGND VPWR _15259_/Q _15063_/Q _10053_/B sky130_fd_sc_hd__nor2_1
X_08909_ VGND VPWR VGND VPWR _15138_/D _15137_/Q _08902_/B _08908_/X _11399_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_66_24 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09889_ VPWR VGND _09970_/A _09893_/A _08862_/C _15477_/D _09024_/A VPWR VGND sky130_fd_sc_hd__o31ai_1
Xhold1240 hold1240/X _14374_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13591__708 VPWR VGND VPWR VGND _14922_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
Xhold1251 hold1251/X _14273_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 _11545_/A _15433_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 _11557_/A _15439_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_745 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1262 hold1262/X _14838_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_1421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11920_ VGND VPWR VGND VPWR _11920_/X _14871_/Q _12229_/A2 _11925_/S _11919_/X sky130_fd_sc_hd__o211a_1
XFILLER_79_1169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11851_ VGND VPWR VGND VPWR _11851_/X _11850_/X _11849_/X _12100_/S _12099_/C1 sky130_fd_sc_hd__a211o_1
Xhold1295 hold1295/X _15285_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_57_1434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10802_ VGND VPWR VPWR VGND _10802_/X _14430_/Q _11216_/S _14686_/Q sky130_fd_sc_hd__mux2_1
X_14570_ _14570_/Q _14570_/CLK _14570_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11782_ VGND VPWR VGND VPWR _11782_/X _11779_/X _11781_/X _12008_/A1 _12017_/C1 sky130_fd_sc_hd__a211o_1
X_13632__749 VPWR VGND VPWR VGND _14972_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_10733_ VPWR VGND VGND VPWR _10733_/X hold466/A _10735_/S sky130_fd_sc_hd__or2_1
XFILLER_18_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10664_ VGND VPWR VPWR VGND _10664_/X hold393/A _10664_/S hold660/A sky130_fd_sc_hd__mux2_1
X_10595_ VPWR VGND VGND VPWR _10595_/X hold335/A _10742_/S sky130_fd_sc_hd__or2_1
X_12403_ VPWR VGND VGND VPWR _12403_/X _14916_/Q _12408_/S sky130_fd_sc_hd__or2_1
X_13485__602 VPWR VGND VPWR VGND _14760_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_15122_ hold837/A _15122_/CLK hold838/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12334_ VGND VPWR VPWR VGND _12334_/X hold826/A _12339_/B hold305/A sky130_fd_sc_hd__mux2_1
XFILLER_31_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13526__643 VPWR VGND VPWR VGND _14806_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_15053_ hold688/A _15053_/CLK _15053_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12265_ VPWR VGND VPWR VGND _12264_/X _12262_/X _12263_/X _12265_/X _12744_/C1 sky130_fd_sc_hd__a22o_1
X_12196_ VPWR VGND VGND VPWR _12177_/Y _12195_/X _10192_/B _15461_/Q _15461_/D _11290_/A
+ sky130_fd_sc_hd__o221a_1
X_11216_ VGND VPWR VPWR VGND _11216_/X _14892_/Q _11216_/S hold463/A sky130_fd_sc_hd__mux2_1
X_11147_ VGND VPWR VGND VPWR _11147_/X hold824/A _11252_/A2 _11146_/X _11143_/S sky130_fd_sc_hd__o211a_1
XFILLER_23_1102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11078_ VGND VPWR VGND VPWR _11078_/X _11075_/X _11077_/X _11252_/C1 _11245_/A1 sky130_fd_sc_hd__a211o_1
X_10029_ VPWR VGND VGND VPWR _10031_/C _10029_/B _15627_/D sky130_fd_sc_hd__nor2_1
X_14906_ hold858/A _14906_/CLK _14906_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14837_ _14837_/Q clkload28/A _14837_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14768_ hold611/A _14768_/CLK _14768_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14699_ hold531/A _14699_/CLK _14699_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07240_ VPWR VGND VGND VPWR _08135_/A _08135_/B _08136_/A sky130_fd_sc_hd__nor2_1
X_07171_ VPWR VGND VGND VPWR _14404_/Q _07301_/A2 _07301_/B1 _07173_/B sky130_fd_sc_hd__o21a_1
X_13269__386 VPWR VGND VPWR VGND _14544_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
Xfanout305 VGND VPWR _10664_/S _10670_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09812_ VGND VPWR VPWR VGND _09830_/S fanout48/X hold1124/X _14240_/D sky130_fd_sc_hd__mux2_2
Xfanout338 VGND VPWR fanout349/X _11261_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout327 VGND VPWR _11146_/B _11142_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout316 VGND VPWR _10972_/S _10994_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout349 VPWR VGND fanout349/X _07893_/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_80_1273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09743_ VGND VPWR VPWR VGND _14303_/D fanout46/X _09760_/S hold246/X sky130_fd_sc_hd__mux2_1
X_09674_ VGND VPWR VPWR VGND _14366_/D hold852/X _09675_/S fanout41/X sky130_fd_sc_hd__mux2_1
XFILLER_76_1309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_08625_ VGND VPWR VGND VPWR _15301_/D hold940/X _08628_/A2 _08624_/X _09977_/A sky130_fd_sc_hd__o211a_1
X_08556_ VPWR VGND VGND VPWR _08605_/A _08977_/B _08556_/Y sky130_fd_sc_hd__nor2_1
X_07507_ VGND VPWR VPWR VGND _15464_/Q _07531_/B _07507_/B sky130_fd_sc_hd__xor2_1
X_08487_ VGND VPWR VGND VPWR _08487_/X hold1336/X _08458_/B _08486_/X _11308_/C1 sky130_fd_sc_hd__o211a_1
X_07438_ VPWR VGND _08548_/B _07507_/B _15459_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_11_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07369_ VPWR VGND VGND VPWR _07369_/X _07369_/A _07369_/B sky130_fd_sc_hd__or2_1
X_13213__330 VPWR VGND VPWR VGND _14488_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
X_09108_ VGND VPWR VPWR VGND _14987_/D hold757/X _09122_/S fanout44/X sky130_fd_sc_hd__mux2_1
X_10380_ VGND VPWR VPWR VGND _10380_/X _14483_/Q _10472_/S hold506/A sky130_fd_sc_hd__mux2_1
X_09039_ VGND VPWR VPWR VGND _15051_/D hold518/X _09053_/S fanout44/X sky130_fd_sc_hd__mux2_1
Xhold381 hold381/X hold381/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 hold370/X hold370/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12050_ VGND VPWR VPWR VGND _12050_/X hold906/A _12220_/S hold820/A sky130_fd_sc_hd__mux2_1
XFILLER_77_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold392 hold392/X hold392/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ VGND VPWR VPWR VGND _11001_/X hold416/A _11231_/S hold542/A sky130_fd_sc_hd__mux2_1
Xfanout861 VGND VPWR _08249_/B2 _07974_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout850 VGND VPWR _10074_/A1 _08278_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout883 VPWR VGND rebuffer7/A _15575_/Q VPWR VGND sky130_fd_sc_hd__buf_6
XFILLER_46_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout872 VGND VPWR _07119_/A _08286_/A VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_13062__179 VPWR VGND VPWR VGND _14305_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
Xhold1081 hold1081/X _14915_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 hold1092/X _14720_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11903_ VGND VPWR VPWR VGND _11903_/X hold773/A _12220_/S hold496/A sky130_fd_sc_hd__mux2_1
Xhold1070 hold1070/X _14350_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_704 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12883_ VPWR VGND VGND VPWR _12883_/A _12883_/B _15604_/D sky130_fd_sc_hd__nor2_1
X_14622_ _14622_/Q _14622_/CLK _14622_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11834_ VPWR VGND VPWR VGND _11833_/X _12175_/A1 _11832_/X _11834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11765_ VPWR VGND VGND VPWR _11765_/X _12098_/A _11765_/B sky130_fd_sc_hd__or2_1
X_14553_ _14553_/Q _14553_/CLK _14553_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_41_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10716_ VPWR VGND VGND VPWR _10716_/X _10732_/S _10716_/B sky130_fd_sc_hd__or2_1
X_14484_ _14484_/Q _14484_/CLK _14484_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11696_ VPWR VGND VGND VPWR _12473_/A _11696_/B _11696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10647_ VGND VPWR VPWR VGND _10647_/X hold645/A _10670_/S hold621/A sky130_fd_sc_hd__mux2_1
Xrebuffer4 VPWR VGND VPWR VGND _07575_/A2 _07486_/C sky130_fd_sc_hd__dlygate4sd1_1
X_10578_ VGND VPWR VPWR VGND _10578_/X _10575_/X _10732_/S _10574_/X sky130_fd_sc_hd__mux2_1
X_15105_ hold904/A _15105_/CLK _15105_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12317_ VGND VPWR VPWR VGND _12317_/X hold970/A _12318_/S hold246/A sky130_fd_sc_hd__mux2_1
X_13760__877 VPWR VGND VPWR VGND _15132_/CLK clkload19/A sky130_fd_sc_hd__inv_2
XFILLER_68_1382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12248_ VGND VPWR VGND VPWR _12248_/X _12245_/X _12247_/X _12580_/A1 _12596_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_29_1322 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15036_ hold555/A _15036_/CLK _15036_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12179_ VGND VPWR VPWR VGND _12179_/X _14363_/Q _12191_/B hold409/A sky130_fd_sc_hd__mux2_1
X_14019__1136 VPWR VGND VPWR VGND _15391_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_9_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_25_907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13654__771 VPWR VGND VPWR VGND _14994_/CLK clkload48/A sky130_fd_sc_hd__inv_2
X_08410_ VGND VPWR VPWR VGND _15367_/D _09658_/A0 _08411_/S hold704/X sky130_fd_sc_hd__mux2_1
X_09390_ VGND VPWR VPWR VGND _14659_/D hold400/X _09411_/S fanout60/X sky130_fd_sc_hd__mux2_1
XFILLER_17_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13948__1065 VPWR VGND VPWR VGND _15320_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_08341_ VGND VPWR VGND VPWR _09556_/C _09240_/A _09311_/B _09198_/C sky130_fd_sc_hd__nand3b_2
X_08272_ VPWR VGND VGND VPWR _08273_/B _14153_/Q _08272_/B sky130_fd_sc_hd__or2_1
X_07223_ VPWR VGND VGND VPWR _12878_/B _07827_/C _10059_/A _07827_/A _07223_/X _15591_/Q
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07154_ VPWR VGND VPWR VGND _07612_/A _07154_/A _07610_/A sky130_fd_sc_hd__or2_2
X_07085_ VPWR VGND VPWR VGND _07769_/A _15545_/Q sky130_fd_sc_hd__inv_2
Xfanout102 VPWR VGND _09825_/A1 _08149_/X VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout113 VGND VPWR _08250_/X _09864_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout146 VGND VPWR _08507_/X _08553_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout135 VPWR VGND VPWR VGND _08726_/C1 _08730_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout124 VGND VPWR _09688_/A0 _08212_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout157 VPWR VGND _09015_/A2 _08936_/X VPWR VGND sky130_fd_sc_hd__buf_2
X_07987_ VGND VPWR VGND VPWR _07987_/X _10072_/B _07985_/X _15081_/Q _07986_/Y sky130_fd_sc_hd__a211o_1
Xfanout168 VGND VPWR _12118_/B1 _12106_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout179 VGND VPWR _12470_/S _12476_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09726_ VGND VPWR VPWR VGND _14317_/D _09726_/A1 _09728_/S hold957/X sky130_fd_sc_hd__mux2_1
X_09657_ VGND VPWR VPWR VGND _14413_/D hold896/X _09657_/S _09691_/A0 sky130_fd_sc_hd__mux2_1
Xtt_um_femto_895 uio_oe[6] tt_um_femto_895/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_76_1139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_09588_ VGND VPWR VPWR VGND _14477_/D hold1027/X _09588_/S _09726_/A1 sky130_fd_sc_hd__mux2_1
X_08608_ VPWR VGND VGND VPWR _07489_/A _08608_/B _08609_/B sky130_fd_sc_hd__nand2b_1
X_08539_ VPWR VGND _15317_/D _08539_/B _08541_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_11550_ VPWR VGND VPWR VGND _11549_/Y _11551_/B _11542_/A _15435_/D sky130_fd_sc_hd__a21oi_1
X_10501_ VGND VPWR VPWR VGND _10501_/X hold631/A _10516_/S hold284/A sky130_fd_sc_hd__mux2_1
X_11481_ VGND VPWR VPWR VGND _11481_/X _15079_/Q _11490_/S _15077_/Q sky130_fd_sc_hd__mux2_1
XFILLER_10_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_12_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10432_ VGND VPWR VPWR VGND _10432_/X hold885/A _10553_/S hold836/A sky130_fd_sc_hd__mux2_1
X_10363_ VPWR VGND VGND VPWR _10363_/X hold411/A _10604_/S sky130_fd_sc_hd__or2_1
X_12102_ VGND VPWR VPWR VGND _12103_/B _12101_/Y _12102_/S _12093_/Y sky130_fd_sc_hd__mux2_1
X_13597__714 VPWR VGND VPWR VGND _14937_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_12033_ VPWR VGND VGND VPWR _12033_/X hold858/A _12112_/S sky130_fd_sc_hd__or2_1
X_10294_ VGND VPWR VPWR VGND _10294_/X hold523/A _10554_/S hold555/A sky130_fd_sc_hd__mux2_1
XFILLER_78_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_667 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_77_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout691 VGND VPWR _08304_/X _08335_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout680 VPWR VGND _09090_/S _09091_/S VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_59_870 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_13638__755 VPWR VGND VPWR VGND _14978_/CLK clkload6/A sky130_fd_sc_hd__inv_2
X_12866_ VGND VPWR VPWR VGND _15590_/D _12866_/A1 _14802_/D _15590_/Q sky130_fd_sc_hd__mux2_1
XFILLER_33_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14605_ hold882/A _14605_/CLK _14605_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11817_ VPWR VGND VGND VPWR _11817_/X hold286/A _12599_/S sky130_fd_sc_hd__or2_1
X_15585_ _15585_/Q clkload43/A _15585_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12797_ VGND VPWR VPWR VGND _12798_/B _08023_/X _12820_/B _08020_/Y sky130_fd_sc_hd__mux2_1
XFILLER_42_781 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_472 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14536_ hold208/A _14536_/CLK _14536_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11748_ VGND VPWR VPWR VGND _11748_/X hold755/A _11748_/S hold511/A sky130_fd_sc_hd__mux2_1
XFILLER_30_998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14467_ hold597/A _14467_/CLK _14467_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11679_ VGND VPWR VPWR VGND _11683_/B hold368/A _12477_/B hold635/A sky130_fd_sc_hd__mux2_1
X_14398_ _14398_/Q clkload54/A _14398_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_08890_ VPWR VGND VGND VPWR _08890_/X _15147_/Q _08918_/B sky130_fd_sc_hd__or2_1
X_15019_ _15019_/Q _15019_/CLK _15019_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07910_ VGND VPWR VGND VPWR _07910_/X _12821_/A _07810_/A _07908_/X _07895_/Y sky130_fd_sc_hd__a211o_2
X_07841_ VGND VPWR _07931_/A _15561_/Q _15562_/Q _07962_/A VPWR VGND sky130_fd_sc_hd__and3_1
X_07772_ VPWR VGND VGND VPWR _07773_/B _15546_/Q _07772_/B sky130_fd_sc_hd__or2_1
XFILLER_42_1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09511_ VGND VPWR VPWR VGND _14548_/D fanout6/X _09513_/S hold455/X sky130_fd_sc_hd__mux2_1
XFILLER_77_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_884 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13390__507 VPWR VGND VPWR VGND _14665_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
X_09442_ VGND VPWR VPWR VGND _14610_/D _09826_/A1 _09449_/S hold462/X sky130_fd_sc_hd__mux2_1
XFILLER_24_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09373_ VGND VPWR VPWR VGND _14673_/D hold397/X _09376_/S _09653_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_75_1172 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14205__923 _14205_/D _14205__923/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_08324_ VGND VPWR VPWR VGND _15495_/D fanout25/X _08338_/S hold917/X sky130_fd_sc_hd__mux2_1
X_13431__548 VPWR VGND VPWR VGND _14706_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_08255_ VPWR VGND VGND VPWR _08214_/A _08094_/X _08254_/X _08255_/X sky130_fd_sc_hd__o21a_1
X_08186_ VGND VPWR _08208_/A _08186_/Y _15549_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07206_ VPWR VGND _07206_/X _07371_/B _15452_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_14_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13284__401 VPWR VGND VPWR VGND _14559_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_07137_ VGND VPWR VGND VPWR _07137_/X _15574_/Q _07141_/A _15572_/Q _12878_/A sky130_fd_sc_hd__or4b_4
XFILLER_58_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13325__442 VPWR VGND VPWR VGND _14600_/CLK clkload41/A sky130_fd_sc_hd__inv_2
XFILLER_60_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_829 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09709_ VGND VPWR VPWR VGND _14334_/D _09710_/S fanout42/X hold1259/X sky130_fd_sc_hd__mux2_4
X_10981_ VGND VPWR VPWR VGND _10981_/X _14211_/Q _10994_/S hold600/A sky130_fd_sc_hd__mux2_1
XFILLER_43_523 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12720_ VGND VPWR VGND VPWR _12720_/X _12720_/A1 _12716_/X _12719_/X _12720_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_15_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12651_ VGND VPWR VPWR VGND _12651_/X _14216_/Q _12651_/S hold171/A sky130_fd_sc_hd__mux2_1
XFILLER_31_729 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11602_ VPWR VGND _11602_/X _11601_/X _11597_/X _12102_/S _11593_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_12582_ VPWR VGND VPWR VGND _12581_/X _12703_/A1 _12580_/X _12582_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_1218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15370_ hold755/A _15370_/CLK _15370_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14018__1135 VPWR VGND VPWR VGND _15390_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_14321_ hold805/A _14321_/CLK _14321_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11533_ VGND VPWR VPWR VGND _11533_/X _11532_/X _11537_/S _15475_/Q sky130_fd_sc_hd__mux2_1
X_11464_ VGND VPWR VPWR VGND _11464_/X _11463_/X _11476_/S _15452_/Q sky130_fd_sc_hd__mux2_1
X_14252_ hold512/A _14252_/CLK _14252_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10415_ VPWR VGND VGND VPWR _10396_/Y _10414_/X _10192_/B _14387_/Q _14387_/D _08735_/C
+ sky130_fd_sc_hd__o221a_1
X_11395_ VPWR VGND VPWR VGND _11392_/B _11368_/A _09938_/A _11395_/X sky130_fd_sc_hd__a21o_1
X_14183_ hold643/A _14183_/CLK _14183_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10346_ VPWR VGND VGND VPWR _10346_/X _10615_/S _10346_/B sky130_fd_sc_hd__or2_1
XFILLER_79_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13947__1064 VPWR VGND VPWR VGND _15319_/CLK clkload26/A sky130_fd_sc_hd__inv_2
X_10277_ VGND VPWR VPWR VGND _10277_/X hold394/A _10602_/S hold240/A sky130_fd_sc_hd__mux2_1
XFILLER_79_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12016_ VPWR VGND VGND VPWR _12016_/X _12106_/S _12016_/B sky130_fd_sc_hd__or2_1
XFILLER_26_1325 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13068__185 VPWR VGND VPWR VGND _14311_/CLK _12972__89/A sky130_fd_sc_hd__inv_2
XFILLER_26_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13872__989 VPWR VGND VPWR VGND _15244_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_15637_ _15637_/Q clkload49/A _15637_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12849_ VGND VPWR VPWR VGND _15573_/D _08236_/X _12860_/S _07141_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15568_ _15568_/Q clkload16/A _15568_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15499_ hold770/A _15499_/CLK _15499_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14519_ hold546/A _14519_/CLK _14519_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13766__883 VPWR VGND VPWR VGND _15138_/CLK _14821_/CLK sky130_fd_sc_hd__inv_2
X_08040_ VPWR VGND VPWR VGND _15619_/Q _08249_/A2 _08051_/B _07426_/X _07331_/A _08039_/X
+ sky130_fd_sc_hd__a221o_1
Xhold903 hold903/X hold903/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 hold925/X hold925/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 hold914/X hold914/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 hold936/X hold936/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 hold947/X hold947/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ VPWR VGND VGND VPWR _09993_/B _09991_/B _15611_/D sky130_fd_sc_hd__nor2_1
Xhold969 hold969/X hold969/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13309__426 VPWR VGND VPWR VGND _14584_/CLK _12957__74/A sky130_fd_sc_hd__inv_2
Xhold958 hold958/X hold958/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08942_ VPWR VGND VPWR VGND _08972_/A hold1447/X _08933_/A _08943_/B _15126_/Q sky130_fd_sc_hd__a22o_1
XFILLER_69_420 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08873_ VGND VPWR VGND VPWR _15156_/D hold1230/X _08893_/A2 _08872_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_07824_ VPWR VGND VPWR VGND _07881_/A2 _07293_/B _10074_/A1 _07824_/X _15088_/Q sky130_fd_sc_hd__a22o_1
XFILLER_77_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07755_ VPWR VGND VPWR VGND _07757_/C _15596_/Q _15549_/Q _07756_/B sky130_fd_sc_hd__a21o_1
XFILLER_77_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_895 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_07686_ _07686_/X _07683_/Y _07684_/X _07685_/X _08249_/B2 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_44_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09425_ VGND VPWR VPWR VGND _14627_/D fanout60/X _09446_/S hold623/X sky130_fd_sc_hd__mux2_1
XFILLER_80_695 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_77_1289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09356_ VGND VPWR VPWR VGND _14690_/D hold991/X _09357_/S clone54/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1418 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08307_ _15512_/D fanout93/X fanout89/X _08305_/Y _08306_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_09287_ VGND VPWR VPWR VGND _14754_/D fanout58/X _09304_/S hold251/X sky130_fd_sc_hd__mux2_1
X_08238_ VGND VPWR VGND VPWR _08250_/B _12214_/A _08172_/X _08237_/X _10058_/A1 sky130_fd_sc_hd__o211a_1
X_08169_ VGND VPWR VGND VPWR _08169_/X _08167_/X _08249_/B2 _08168_/X sky130_fd_sc_hd__a21bo_1
X_10200_ VGND VPWR VPWR VGND _10200_/X _10197_/X _10995_/S _10196_/X sky130_fd_sc_hd__mux2_1
X_11180_ VGND VPWR VGND VPWR _11180_/X _11179_/X _11178_/X _11170_/S _11180_/C1 sky130_fd_sc_hd__a211o_1
X_10131_ VGND VPWR VPWR VGND _10131_/X hold520/A _10353_/S hold309/A sky130_fd_sc_hd__mux2_1
X_10062_ VPWR VGND VPWR VGND _10062_/B _10062_/D _10062_/C _10062_/A _10063_/D sky130_fd_sc_hd__or4_1
X_14870_ hold910/A _14870_/CLK _14870_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13102__219 VPWR VGND VPWR VGND _14345_/CLK _12970__87/A sky130_fd_sc_hd__inv_2
XFILLER_56_1329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12703_ VGND VPWR VGND VPWR _12703_/X _12703_/A1 _12698_/X _12702_/X _12864_/A1 sky130_fd_sc_hd__o211a_1
X_10964_ VGND VPWR VPWR VGND _10964_/X hold772/A _10964_/S hold346/A sky130_fd_sc_hd__mux2_1
X_10895_ VPWR VGND VGND VPWR _10895_/X _14400_/Q _12380_/B sky130_fd_sc_hd__or2_1
X_13453__570 VPWR VGND VPWR VGND _14728_/CLK clkload40/A sky130_fd_sc_hd__inv_2
X_12634_ VGND VPWR VPWR VGND _12634_/X hold824/A _12635_/B hold421/A sky130_fd_sc_hd__mux2_1
X_15422_ hold711/A _15422_/CLK _15422_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15353_ _15353_/Q _15353_/CLK _15353_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12565_ VPWR VGND VPWR VGND _12564_/X _12658_/A _12713_/B1 _12565_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_773 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14304_ _14304_/Q _14304_/CLK _14304_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11516_ VGND VPWR VPWR VGND _15089_/D _11515_/X _11528_/S hold1426/X sky130_fd_sc_hd__mux2_1
XFILLER_32_1373 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15284_ _15284_/Q _15284_/CLK _15284_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12496_ VGND VPWR VPWR VGND _12496_/X hold740/A _12652_/S hold467/A sky130_fd_sc_hd__mux2_1
XFILLER_50_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14235_ hold185/A _14235_/CLK _14235_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11447_ VGND VPWR VPWR VGND _15066_/D _11446_/X _11477_/S hold1415/X sky130_fd_sc_hd__mux2_1
X_11378_ VGND VPWR VPWR VGND _11378_/X _11377_/X _11387_/S _14847_/Q sky130_fd_sc_hd__mux2_1
X_13800__917 VPWR VGND VPWR VGND _15172_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_14166_ hold651/A _14166_/CLK _14166_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10329_ VGND VPWR VPWR VGND _10333_/B hold797/A _11102_/S hold495/A sky130_fd_sc_hd__mux2_1
XFILLER_79_773 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07540_ VGND VPWR VGND VPWR _07539_/Y _07523_/Y _07518_/X _07552_/B1 _07560_/B _15565_/Q
+ sky130_fd_sc_hd__a32oi_4
XFILLER_47_692 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_35_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14999_ _14999_/Q _14999_/CLK _14999_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07471_ VPWR VGND VGND VPWR _15448_/Q _07471_/B _07486_/B sky130_fd_sc_hd__nor2_1
X_09210_ VGND VPWR VPWR VGND _14883_/D hold769/X _09228_/S fanout50/X sky130_fd_sc_hd__mux2_1
X_09141_ VGND VPWR VPWR VGND _14957_/D fanout54/X _09157_/S hold831/X sky130_fd_sc_hd__mux2_1
X_09072_ VGND VPWR VPWR VGND _15021_/D hold1095/X _09090_/S fanout54/X sky130_fd_sc_hd__mux2_1
X_08023_ VPWR VGND VGND VPWR _08023_/X _08023_/A _08023_/B sky130_fd_sc_hd__or2_1
XFILLER_11_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold700 hold700/X hold700/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold711 hold711/X hold711/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 hold733/X hold733/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 hold744/X hold744/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 hold722/X hold722/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 hold755/X hold755/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 hold766/X hold766/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 hold777/X hold777/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 hold788/X hold788/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ VPWR VGND VGND VPWR _15478_/D _09974_/A _09974_/B sky130_fd_sc_hd__or2_1
Xhold799 hold799/X hold799/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08925_ VGND VPWR VGND VPWR _15130_/D _15129_/Q _08902_/B _08924_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
Xhold1400 hold1400/X _14893_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14017__1134 VPWR VGND VPWR VGND _15389_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_08856_ VPWR VGND VGND VPWR _08859_/C _14146_/Q hold149/A sky130_fd_sc_hd__or2_1
Xhold1433 _09234_/A _14808_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 hold1411/X _15145_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold1422 hold1422/X _15092_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13396__513 VPWR VGND VPWR VGND _14671_/CLK clkload34/A sky130_fd_sc_hd__inv_2
Xhold1444 hold1444/X _15321_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _08468_/A _15342_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1466 _08920_/A _15132_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07807_ VGND VPWR VPWR VGND _07808_/B _15593_/Q _07807_/S _07519_/B sky130_fd_sc_hd__mux2_1
X_08787_ VGND VPWR VPWR VGND _15222_/D _08808_/S clone47/A hold1164/X sky130_fd_sc_hd__mux2_4
X_07738_ VPWR VGND _07738_/X _07739_/B _15555_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_13437__554 VPWR VGND VPWR VGND _14712_/CLK clkload18/A sky130_fd_sc_hd__inv_2
XFILLER_53_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07669_ VGND VPWR VPWR VGND _07669_/X _15091_/Q _07881_/A2 _07339_/B _07972_/B sky130_fd_sc_hd__o2bb2a_1
X_09408_ VGND VPWR VPWR VGND _14641_/D hold606/X _09408_/S _09827_/A1 sky130_fd_sc_hd__mux2_1
X_10680_ VGND VPWR VPWR VGND _10680_/X hold613/A _10687_/B hold442/A sky130_fd_sc_hd__mux2_1
XFILLER_13_548 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13946__1063 VPWR VGND VPWR VGND _15318_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_09339_ VGND VPWR VPWR VGND _14705_/D hold491/X _09342_/S _09653_/A0 sky130_fd_sc_hd__mux2_1
X_12350_ VGND VPWR VGND VPWR _12350_/X hold973/A _12861_/A1 _12375_/S _12349_/X sky130_fd_sc_hd__o211a_1
X_11301_ VPWR VGND _11307_/B _11302_/B _11302_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_12281_ VGND VPWR VPWR VGND _12281_/X _14206_/Q _12282_/S hold172/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11232_ VGND VPWR VPWR VGND _11232_/X _14346_/Q _11240_/S _15258_/Q sky130_fd_sc_hd__mux2_1
XFILLER_20_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11163_ VPWR VGND VPWR VGND _11162_/X _11181_/A1 _11161_/X _11163_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10114_ VPWR VGND VGND VPWR _10114_/X hold532/A _10609_/S sky130_fd_sc_hd__or2_1
X_11094_ VPWR VGND VGND VPWR _11094_/X _14310_/Q _11107_/S sky130_fd_sc_hd__or2_1
XFILLER_62_1344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10045_ VGND VPWR _10049_/B _15635_/Q _15634_/Q _10045_/C VPWR VGND sky130_fd_sc_hd__and3_1
X_14922_ hold540/A _14922_/CLK _14922_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14853_ _14853_/Q clkload26/A _14853_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_1041 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14784_ hold608/A _14784_/CLK _14784_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11996_ VPWR VGND VGND VPWR _11996_/X hold322/A _12006_/B sky130_fd_sc_hd__or2_1
XFILLER_16_342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10947_ VGND VPWR VGND VPWR _10947_/X _11178_/C1 _10943_/X _10946_/X _11180_/C1 sky130_fd_sc_hd__o211a_1
X_10878_ VPWR VGND VPWR VGND _10877_/X _10333_/A _10891_/C1 _10878_/X sky130_fd_sc_hd__a21o_1
X_15405_ hold818/A _15405_/CLK _15405_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12617_ VGND VPWR VGND VPWR _12617_/X _12737_/B1 _12613_/X _12616_/X _12739_/C1 sky130_fd_sc_hd__o211a_1
X_15336_ _15336_/Q _15336_/CLK _15336_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12548_ VPWR VGND VGND VPWR _12548_/X hold310/A _12664_/S sky130_fd_sc_hd__or2_1
X_15267_ _15267_/Q _15267_/CLK _15267_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 _07593_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_13230__347 VPWR VGND VPWR VGND _14505_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_12479_ VGND VPWR VPWR VGND _12479_/X hold964/A _12479_/S hold711/A sky130_fd_sc_hd__mux2_1
XFILLER_67_1200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14218_ _14218_/Q _14218_/CLK _14218_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15198_ hold190/A _15198_/CLK _15198_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14149_ hold226/A _14149_/CLK _14149_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout509 VPWR VGND _12716_/S fanout539/X VPWR VGND sky130_fd_sc_hd__buf_2
X_13878__995 VPWR VGND VPWR VGND _15250_/CLK clkload42/A sky130_fd_sc_hd__inv_2
X_13083__200 VPWR VGND VPWR VGND _14326_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_08710_ VGND VPWR VGND VPWR _15278_/D hold1036/X _08721_/A2 _08709_/X _11294_/A sky130_fd_sc_hd__o211a_1
X_09690_ VGND VPWR VPWR VGND _14350_/D hold1070/X _09690_/S _09690_/A0 sky130_fd_sc_hd__mux2_1
X_13124__241 VPWR VGND VPWR VGND _14367_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_08641_ VPWR VGND VGND VPWR _08640_/X _08690_/S _08194_/Y _14408_/Q _08641_/X _08639_/X
+ sky130_fd_sc_hd__o221a_1
Xrebuffer14 VPWR VGND VPWR VGND _07564_/B _07479_/Y sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer25 VPWR VGND VPWR VGND rebuffer25/X rebuffer26/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer36 VPWR VGND VPWR VGND rebuffer36/X rebuffer37/X sky130_fd_sc_hd__dlygate4sd1_1
X_08572_ VPWR VGND VPWR VGND _15598_/Q _15453_/Q _07494_/X _08586_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07523_ VPWR VGND VGND VPWR _07523_/Y _07523_/B _07534_/A sky130_fd_sc_hd__nor2_4
X_07454_ VGND VPWR VGND VPWR _07454_/X _15454_/Q _15599_/Q _07496_/A _07453_/X sky130_fd_sc_hd__o211a_1
XFILLER_62_481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07385_ VPWR VGND VGND VPWR _07971_/A _07385_/Y _07981_/A sky130_fd_sc_hd__nand2_1
X_09124_ VGND VPWR VPWR VGND _14971_/D hold327/X _09124_/S _09689_/A0 sky130_fd_sc_hd__mux2_1
X_09055_ VGND VPWR VPWR VGND _15035_/D hold768/X _09055_/S _09655_/A0 sky130_fd_sc_hd__mux2_1
X_12988__105 VPWR VGND VPWR VGND _14231_/CLK clkload20/A sky130_fd_sc_hd__inv_2
X_08006_ VPWR VGND VPWR VGND _08006_/B _08006_/C _08010_/A _08007_/B sky130_fd_sc_hd__or3_1
XFILLER_11_1265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold530 hold530/X hold530/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 hold541/X hold541/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 hold563/X hold563/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_739 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold552 hold552/X hold552/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 hold596/X hold596/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 hold585/X hold585/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 hold574/X hold574/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ VPWR VGND VGND VPWR hold1274/X _09937_/B _08529_/A _14766_/D sky130_fd_sc_hd__o21a_1
X_08908_ VPWR VGND VGND VPWR _08908_/X _15138_/Q _08924_/B sky130_fd_sc_hd__or2_1
X_09888_ VGND VPWR VPWR VGND _14147_/D hold1228/X _09888_/S _09887_/X sky130_fd_sc_hd__mux2_1
Xhold1230 hold1230/X _15155_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 hold1241/X _15134_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 hold1252/X _14311_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 _11563_/A _15442_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 hold1274/X _14763_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1263 hold1263/X _14304_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_990 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08839_ VGND VPWR VPWR VGND _15174_/D fanout14/X _08850_/S hold367/X sky130_fd_sc_hd__mux2_1
Xhold1296 hold1296/X _14846_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11850_ VGND VPWR VPWR VGND _11850_/X hold827/A _12089_/S hold818/A sky130_fd_sc_hd__mux2_1
X_10801_ VGND VPWR VGND VPWR _10801_/X _11217_/C1 _10796_/X _10800_/X _10765_/S sky130_fd_sc_hd__o211a_1
X_13671__788 VPWR VGND VPWR VGND _15011_/CLK clkload14/A sky130_fd_sc_hd__inv_2
X_11781_ VGND VPWR VGND VPWR _11781_/X hold958/A _12188_/A2 _11995_/S _11780_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10732_ VGND VPWR VPWR VGND _10732_/X _10731_/X _10732_/S _10730_/X sky130_fd_sc_hd__mux2_1
X_10663_ VGND VPWR VGND VPWR _10663_/X _10667_/C1 _10662_/X _10659_/X _10737_/C1 sky130_fd_sc_hd__o211a_1
X_12402_ VGND VPWR VPWR VGND _12402_/X _12401_/X _12721_/S _12400_/X sky130_fd_sc_hd__mux2_1
X_10594_ VGND VPWR VPWR VGND _10594_/X hold372/A _10742_/S hold701/A sky130_fd_sc_hd__mux2_1
X_15121_ _15121_/Q _15121_/CLK _15121_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12333_ VGND VPWR VGND VPWR _12333_/X _12596_/C1 _12328_/X _12332_/X _12740_/C1 sky130_fd_sc_hd__o211a_1
X_13565__682 VPWR VGND VPWR VGND _14896_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_15052_ hold707/A _15052_/CLK _15052_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_3_0_clk clkload1/A clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_12264_ VGND VPWR VPWR VGND _12264_/X _12261_/X _12328_/S _12260_/X sky130_fd_sc_hd__mux2_1
X_11215_ VGND VPWR VGND VPWR _11215_/X hold932/A _11215_/A2 _11214_/X _11215_/C1 sky130_fd_sc_hd__o211a_1
X_12195_ VPWR VGND VPWR VGND _12194_/X _12029_/A _12195_/B1 _12195_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_11146_ VPWR VGND VGND VPWR _11146_/X hold421/A _11146_/B sky130_fd_sc_hd__or2_1
XFILLER_49_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11077_ VGND VPWR VGND VPWR _11077_/X _15025_/Q _11252_/A2 _11076_/X _11250_/S sky130_fd_sc_hd__o211a_1
X_13108__225 VPWR VGND VPWR VGND _14351_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_10028_ VPWR VGND VGND VPWR _10028_/A _10028_/B _10029_/B sky130_fd_sc_hd__nor2_1
X_14905_ hold322/A _14905_/CLK _14905_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14836_ _14836_/Q clkload28/A _14836_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14767_ _14767_/Q _14767_/CLK _14767_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11979_ VPWR VGND VGND VPWR _11979_/X _12106_/S _11979_/B sky130_fd_sc_hd__or2_1
X_14698_ _14698_/Q _14698_/CLK _14698_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_07170_ VPWR VGND VPWR VGND _07668_/A _07167_/Y _07338_/A _07170_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_197 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14016__1133 VPWR VGND VPWR VGND _15388_/CLK clkload36/A sky130_fd_sc_hd__inv_2
X_15319_ _15319_/Q _15319_/CLK _15319_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13806__923 VPWR VGND VPWR VGND _15178_/CLK clkload17/A sky130_fd_sc_hd__inv_2
Xfanout339 VPWR VGND _11223_/S fanout349/X VPWR VGND sky130_fd_sc_hd__buf_2
X_09811_ VGND VPWR VPWR VGND _14241_/D _09827_/S clone46/X hold1140/X sky130_fd_sc_hd__mux2_4
Xfanout306 VGND VPWR _10664_/S _10720_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout328 VGND VPWR _10964_/S _11146_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout317 VPWR VGND _10972_/S _11231_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_13945__1062 VPWR VGND VPWR VGND _15317_/CLK clkload28/A sky130_fd_sc_hd__inv_2
X_09742_ VGND VPWR VPWR VGND _14304_/D _09760_/S fanout48/X hold1263/X sky130_fd_sc_hd__mux2_4
XFILLER_80_1285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_41_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09673_ VGND VPWR VPWR VGND _14367_/D hold880/X _09687_/S fanout45/X sky130_fd_sc_hd__mux2_1
X_08624_ VGND VPWR VGND VPWR _08624_/X _08626_/A _08627_/C1 hold960/X _08623_/Y sky130_fd_sc_hd__a211o_1
X_08555_ VGND VPWR VPWR VGND _08977_/B _15557_/Q _08591_/B _08604_/B2 _08554_/Y sky130_fd_sc_hd__o2bb2a_1
X_07506_ VPWR VGND VGND VPWR _07506_/A _07530_/B _07545_/A sky130_fd_sc_hd__nor2_1
X_08486_ VPWR VGND VGND VPWR _08486_/X _15333_/Q _08486_/B sky130_fd_sc_hd__or2_1
X_07437_ VGND VPWR _07507_/B _08548_/A _15460_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07368_ VPWR VGND VGND VPWR _08201_/B _07368_/A _12845_/A sky130_fd_sc_hd__or2_1
X_13549__666 VPWR VGND VPWR VGND _14880_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_09107_ VGND VPWR VPWR VGND _14988_/D hold748/X _09124_/S clone100/X sky130_fd_sc_hd__mux2_1
X_07299_ VGND VPWR _07301_/A2 _07301_/B1 _07300_/B _14400_/Q VPWR VGND sky130_fd_sc_hd__o21ai_1
X_09038_ VGND VPWR VPWR VGND _15052_/D hold707/X _09055_/S clone100/X sky130_fd_sc_hd__mux2_1
Xhold371 hold371/X hold371/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_536 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold360 hold360/X hold360/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 hold393/X hold393/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 hold382/X hold382/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ VGND VPWR VGND VPWR _11000_/X _10997_/X _10999_/X _11004_/A1 _11235_/C1 sky130_fd_sc_hd__a211o_1
Xfanout840 VPWR VGND _07544_/B fanout844/X VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_77_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xfanout851 VGND VPWR _07417_/X _10074_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout884 VPWR VGND _07765_/B _07141_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout862 VGND VPWR _07136_/Y _08249_/B2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout873 VPWR VGND _07331_/A _15583_/Q VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_46_713 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1060 hold1060/X _15505_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ VPWR VGND VPWR VGND _08233_/B _08073_/B _08198_/S _12883_/B sky130_fd_sc_hd__a21oi_1
XFILLER_45_234 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1071 hold1071/X _15507_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 hold1093/X _15023_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ VGND VPWR VPWR VGND _11902_/X _14484_/Q _12220_/S hold453/A sky130_fd_sc_hd__mux2_1
Xhold1082 hold1082/X _15016_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14621_ hold619/A _14621_/CLK _14621_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11833_ VGND VPWR VPWR VGND _11833_/X _11830_/X _12174_/S _11829_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_1274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14552_ hold640/A _14552_/CLK _14552_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11764_ VGND VPWR VPWR VGND _11764_/X hold434/A _12086_/S hold390/A sky130_fd_sc_hd__mux2_1
XFILLER_13_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14483_ _14483_/Q _14483_/CLK _14483_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10715_ VGND VPWR VPWR VGND _10715_/X hold584/A _10743_/B hold237/A sky130_fd_sc_hd__mux2_1
X_11695_ VGND VPWR VPWR VGND _11696_/B _11694_/Y _12472_/S _11686_/Y sky130_fd_sc_hd__mux2_1
XFILLER_9_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_14_687 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_70_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12979__96 VPWR VGND VPWR VGND _14222_/CLK _12979__96/A sky130_fd_sc_hd__inv_2
X_10646_ VGND VPWR VPWR VGND _10650_/B hold721/A _10670_/S hold159/A sky130_fd_sc_hd__mux2_1
X_15104_ _15104_/Q _15104_/CLK _15104_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10577_ VGND VPWR VGND VPWR _10577_/X _10745_/A1 _10573_/X _10576_/X _10741_/C1 sky130_fd_sc_hd__o211a_1
X_12316_ VGND VPWR VPWR VGND _12320_/B hold706/A _12318_/S hold244/A sky130_fd_sc_hd__mux2_1
X_12247_ VGND VPWR VGND VPWR _12247_/X hold908/A _12705_/A2 _12581_/S _12246_/X sky130_fd_sc_hd__o211a_1
X_15035_ hold768/A _15035_/CLK _15035_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_69_849 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12178_ VGND VPWR VPWR VGND _12178_/X hold998/A _12191_/B hold536/A sky130_fd_sc_hd__mux2_1
X_13342__459 VPWR VGND VPWR VGND _14617_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
X_11129_ VGND VPWR VPWR VGND _11129_/X _14215_/Q _11146_/B _15223_/Q sky130_fd_sc_hd__mux2_1
XFILLER_37_757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13195__312 VPWR VGND VPWR VGND _14470_/CLK clkload51/A sky130_fd_sc_hd__inv_2
X_14819_ _14819_/Q _14821_/CLK _14819_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_08340_ VPWR VGND VGND VPWR _15639_/Q _09729_/A _09834_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_974 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_71_1229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08271_ VGND VPWR _08113_/X _08270_/X _08271_/Y _08214_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
X_13236__353 VPWR VGND VPWR VGND _14511_/CLK clkload35/A sky130_fd_sc_hd__inv_2
X_07222_ VGND VPWR VGND VPWR _10061_/A _07222_/B _07222_/A sky130_fd_sc_hd__xnor2_4
X_07153_ VPWR VGND VGND VPWR _15475_/Q _07153_/B _07610_/A sky130_fd_sc_hd__nor2_1
X_07084_ VPWR VGND VPWR VGND _07736_/A _15556_/Q sky130_fd_sc_hd__inv_2
Xfanout103 VPWR VGND VPWR VGND _09859_/A0 _08149_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout136 VPWR VGND _08534_/B1 _08540_/B1 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout125 VGND VPWR _08190_/X _09792_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout147 VGND VPWR _08686_/A2 _08701_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout114 VGND VPWR _09622_/A1 _08250_/X VPWR VGND sky130_fd_sc_hd__buf_1
Xfanout158 VGND VPWR _11421_/X _11431_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_07986_ VPWR VGND VGND VPWR _07981_/A _10075_/A _07984_/X _07333_/Y _07986_/Y sky130_fd_sc_hd__o22ai_1
Xfanout169 VGND VPWR _08298_/A1 _12118_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09725_ VGND VPWR VPWR VGND _14318_/D _09864_/A0 _09725_/S hold476/X sky130_fd_sc_hd__mux2_1
XFILLER_55_543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09656_ VGND VPWR VPWR VGND _14414_/D hold833/X _09656_/S _09690_/A0 sky130_fd_sc_hd__mux2_1
X_08607_ VGND VPWR VGND VPWR _15306_/D hold1052/X _08613_/A2 _08606_/X _11337_/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xtt_um_femto_896 uio_oe[7] tt_um_femto_896/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_09587_ VGND VPWR VPWR VGND _14478_/D hold863/X _09587_/S _09864_/A0 sky130_fd_sc_hd__mux2_1
X_08538_ VPWR VGND VPWR VGND _08540_/B1 _15316_/Q _08540_/A2 _08539_/B hold1414/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_248 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08469_ VGND VPWR VGND VPWR _15342_/D hold1162/X _08483_/A2 _08468_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_10500_ VGND VPWR VPWR VGND _10500_/X _14198_/Q _10516_/S hold341/A sky130_fd_sc_hd__mux2_1
X_11480_ VGND VPWR VPWR VGND _15077_/D _11479_/X _11480_/S _15077_/Q sky130_fd_sc_hd__mux2_1
X_10431_ VGND VPWR VGND VPWR _10431_/X _10717_/C1 _10426_/X _10430_/X clone2/X sky130_fd_sc_hd__o211a_1
X_10362_ VGND VPWR VPWR VGND _10362_/X _10361_/X _10625_/S _10360_/X sky130_fd_sc_hd__mux2_1
X_10293_ VGND VPWR VGND VPWR _10293_/X _10634_/C1 _10288_/X _10292_/X _10626_/C1 sky130_fd_sc_hd__o211a_1
X_12101_ VPWR VGND VPWR VGND _12100_/X _12101_/A1 _12099_/X _12101_/Y sky130_fd_sc_hd__a21oi_1
X_12032_ VGND VPWR VPWR VGND _12032_/X _12031_/X _12106_/S _12030_/X sky130_fd_sc_hd__mux2_1
Xhold190 hold190/X hold190/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout692 VPWR VGND _08902_/B _08880_/B VPWR VGND sky130_fd_sc_hd__buf_2
X_14015__1132 VPWR VGND VPWR VGND _15387_/CLK clkload45/A sky130_fd_sc_hd__inv_2
Xfanout681 VPWR VGND _09088_/S _09091_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_13677__794 VPWR VGND VPWR VGND _15017_/CLK clkload55/A sky130_fd_sc_hd__inv_2
Xfanout670 VPWR VGND _09188_/S _09164_/X VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_74_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12865_ VGND VPWR VPWR VGND _15589_/D _12584_/A _12870_/S _15589_/Q sky130_fd_sc_hd__mux2_1
XFILLER_61_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11816_ VGND VPWR VPWR VGND _11816_/X hold398/A _12589_/S hold235/A sky130_fd_sc_hd__mux2_1
X_12796_ VPWR VGND _15556_/D _09976_/B _15556_/Q _09975_/A _12795_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_15584_ VGND VPWR VGND VPWR _15584_/Q _15584_/D clkload27/A sky130_fd_sc_hd__dfxtp_4
X_14604_ hold519/A _14604_/CLK _14604_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_30_900 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14535_ hold421/A _14535_/CLK _14535_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11747_ VGND VPWR VGND VPWR _11747_/X _15485_/Q _12861_/A1 _12396_/S _11746_/X sky130_fd_sc_hd__o211a_1
X_13944__1061 VPWR VGND VPWR VGND _15316_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_11678_ VPWR VGND VGND VPWR _11659_/Y _11677_/X _10192_/B _15447_/Q _15447_/D _11420_/S
+ sky130_fd_sc_hd__o221a_1
X_14466_ hold716/A _14466_/CLK _14466_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14397_ _14397_/Q clkload53/A _14397_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_10629_ VGND VPWR VGND VPWR _10629_/X hold917/A _10629_/A2 _10628_/X _10625_/S sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15018_ _15018_/Q _15018_/CLK _15018_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07840_ VPWR VGND _07962_/A _07990_/A _15560_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07771_ VPWR VGND _08247_/A _07770_/B _08272_/B _14153_/Q _07766_/Y VGND VPWR sky130_fd_sc_hd__a31o_1
X_09510_ VGND VPWR VPWR VGND _14549_/D fanout9/X _09520_/S hold877/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_1397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_37_554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_77_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09441_ VGND VPWR VPWR VGND _14611_/D _09825_/A1 _09441_/S hold806/X sky130_fd_sc_hd__mux2_1
XFILLER_24_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09372_ VGND VPWR VPWR VGND _14674_/D hold435/X _09379_/S _09548_/A1 sky130_fd_sc_hd__mux2_1
X_08323_ VGND VPWR VPWR VGND _15496_/D fanout28/X _08338_/S hold936/X sky130_fd_sc_hd__mux2_1
X_13470__587 VPWR VGND VPWR VGND _14745_/CLK clkload8/A sky130_fd_sc_hd__inv_2
X_08254_ VPWR VGND VGND VPWR _08173_/Y _08253_/X _08172_/X _12222_/C1 _08254_/X _10058_/A1
+ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07205_ VGND VPWR VPWR VGND _07220_/S _15597_/Q _14386_/Q _07371_/B sky130_fd_sc_hd__mux2_2
X_08185_ VPWR VGND VPWR VGND _08182_/X _08280_/B2 _08184_/X _08185_/Y sky130_fd_sc_hd__a21oi_1
X_07136_ VPWR VGND VGND VPWR _15574_/Q _12878_/A _07136_/Y _15572_/Q _07141_/A sky130_fd_sc_hd__nor4b_1
X_13364__481 VPWR VGND VPWR VGND _14639_/CLK clkload34/A sky130_fd_sc_hd__inv_2
XFILLER_48_808 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09708_ VGND VPWR VPWR VGND _14335_/D fanout46/X _09710_/S hold829/X sky130_fd_sc_hd__mux2_1
XFILLER_60_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07969_ VPWR VGND VPWR VGND _10064_/A _07942_/C _07345_/X _07983_/A _07968_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_21_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10980_ VGND VPWR VPWR VGND _10980_/X hold507/A _10994_/S hold293/A sky130_fd_sc_hd__mux2_1
X_09639_ VGND VPWR VPWR VGND _14431_/D hold785/X _09656_/S fanout45/X sky130_fd_sc_hd__mux2_1
X_13711__828 VPWR VGND VPWR VGND _15051_/CLK clkload51/A sky130_fd_sc_hd__inv_2
XFILLER_43_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12650_ VGND VPWR VPWR VGND _12650_/X hold535/A _12652_/S hold262/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11601_ VGND VPWR VGND VPWR _11601_/X _11598_/X _11600_/X _11995_/S _12017_/C1 sky130_fd_sc_hd__a211o_1
X_12581_ VGND VPWR VPWR VGND _12581_/X _12578_/X _12581_/S _12577_/X sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14320_ hold689/A _14320_/CLK _14320_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11532_ VGND VPWR VPWR VGND _11532_/X _15096_/Q _11535_/C _15094_/Q sky130_fd_sc_hd__mux2_1
X_12949__66 VPWR VGND VPWR VGND _14192_/CLK _12981__98/A sky130_fd_sc_hd__inv_2
XFILLER_23_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11463_ VGND VPWR VPWR VGND _11463_/X _15073_/Q _11475_/S _15071_/Q sky130_fd_sc_hd__mux2_1
X_14251_ hold366/A _14251_/CLK _14251_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14182_ _14182_/Q _14182_/CLK _14182_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10414_ VPWR VGND VPWR VGND _10413_/X _10507_/A _12195_/B1 _10414_/X sky130_fd_sc_hd__a21o_1
X_11394_ VGND VPWR VPWR VGND _14851_/D _11393_/X _11398_/A _14851_/Q sky130_fd_sc_hd__mux2_1
X_13605__722 VPWR VGND VPWR VGND _14945_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_10345_ VGND VPWR VPWR VGND _10345_/X hold665/A _10687_/B hold173/A sky130_fd_sc_hd__mux2_1
XFILLER_79_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10276_ VGND VPWR VPWR VGND _10280_/B hold534/A _10602_/S hold229/A sky130_fd_sc_hd__mux2_1
XFILLER_79_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12015_ VGND VPWR VPWR VGND _12015_/X hold735/A _12112_/S hold307/A sky130_fd_sc_hd__mux2_1
XFILLER_2_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_6_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_14187__905 _14187_/D _14187__905/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_46_351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12848_ VGND VPWR VPWR VGND _15572_/D _08253_/X _12860_/S _15572_/Q sky130_fd_sc_hd__mux2_1
X_15636_ _15636_/Q clkload49/A _15636_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12779_ VGND VPWR _12777_/X _12778_/X _12779_/Y _12776_/Y VPWR VGND sky130_fd_sc_hd__o21ai_1
X_15567_ _15567_/Q clkload16/A _15567_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_9_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14518_ hold236/A _14518_/CLK _14518_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15498_ hold926/A _15498_/CLK _15498_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14449_ hold862/A _14449_/CLK _14449_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold904 hold904/X hold904/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold915 hold915/X hold915/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 hold937/X hold937/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 hold926/X hold926/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13348__465 VPWR VGND VPWR VGND _14623_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
Xhold948 hold948/X hold948/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12963__80 VPWR VGND VPWR VGND _14206_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_09990_ VPWR VGND VPWR VGND _09989_/C _15610_/Q hold1320/X _09991_/B sky130_fd_sc_hd__a21oi_1
Xhold959 hold959/X hold959/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08941_ VPWR VGND _15127_/D _08941_/B _08955_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08872_ VPWR VGND VGND VPWR _08872_/X _08872_/A _08918_/B sky130_fd_sc_hd__or2_1
X_07823_ VGND VPWR VGND VPWR _07668_/B _07820_/A _07859_/B _07823_/X _07291_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07754_ VGND VPWR _07754_/X _15596_/Q _15549_/Q _07757_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_77_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_682 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_811 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07685_ VGND VPWR VGND VPWR _10074_/A1 _07679_/A _07859_/B _07685_/X _07174_/Y sky130_fd_sc_hd__a2bb2o_1
XFILLER_77_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09424_ VGND VPWR VPWR VGND _14628_/D fanout65/X _09443_/S hold579/X sky130_fd_sc_hd__mux2_1
XFILLER_52_365 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09355_ VGND VPWR VPWR VGND _14691_/D hold754/X _09376_/S fanout60/X sky130_fd_sc_hd__mux2_1
X_08306_ VPWR VGND VGND VPWR _08306_/X _08306_/A _08318_/S sky130_fd_sc_hd__or2_1
X_09286_ VGND VPWR VPWR VGND _14755_/D fanout60/X _09307_/S hold413/X sky130_fd_sc_hd__mux2_1
X_08237_ VPWR VGND VGND VPWR _08173_/Y _08234_/X _08198_/S _08236_/X _08237_/X sky130_fd_sc_hd__o22a_1
X_14014__1131 VPWR VGND VPWR VGND _15386_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_08168_ VPWR VGND VGND VPWR _07886_/A _08153_/X _08147_/A _08155_/X _08168_/X sky130_fd_sc_hd__o22a_1
XFILLER_69_36 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_08099_ VGND VPWR _08099_/B _08099_/Y _15553_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07119_ VPWR VGND VPWR VGND _07119_/Y _07119_/A sky130_fd_sc_hd__inv_2
X_10130_ VGND VPWR VPWR VGND _10130_/X _14188_/Q _10612_/S hold186/A sky130_fd_sc_hd__mux2_1
X_10061_ VPWR VGND VPWR VGND _10061_/B _10061_/D _10061_/C _10061_/A _10062_/D sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_8_Left_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13943__1060 VPWR VGND VPWR VGND _15315_/CLK clkload29/A sky130_fd_sc_hd__inv_2
XFILLER_76_958 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_60_1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13141__258 VPWR VGND VPWR VGND _14416_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_10963_ VGND VPWR VGND VPWR _10963_/X _10960_/X _10962_/X _11178_/C1 _11180_/C1 sky130_fd_sc_hd__a211o_1
X_12702_ VGND VPWR VGND VPWR _12702_/X _12701_/X _12700_/X _12698_/S _12702_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_16_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10894_ VPWR VGND VPWR VGND _10894_/X _11210_/A _10867_/X _10875_/X _10893_/X _10892_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_31_527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15421_ hold425/A _15421_/CLK _15421_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_16_579 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12633_ VGND VPWR VGND VPWR _12633_/X _12630_/X _12632_/X _12737_/B1 _12740_/A1 sky130_fd_sc_hd__a211o_1
X_15352_ _15352_/Q _15352_/CLK _15352_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12564_ VPWR VGND _12564_/X _12563_/X _12559_/X _12694_/S _12555_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_15_1027 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14303_ hold246/A _14303_/CLK _14303_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11515_ VGND VPWR VPWR VGND _11515_/X _11514_/X _11530_/S _15469_/Q sky130_fd_sc_hd__mux2_1
X_15283_ hold953/A _15283_/CLK _15283_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_11_262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13035__152 VPWR VGND VPWR VGND _14278_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_14234_ hold159/A _14234_/CLK _14234_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12495_ VGND VPWR VPWR VGND _12495_/X hold662/A _12652_/S hold289/A sky130_fd_sc_hd__mux2_1
X_11446_ VGND VPWR VPWR VGND _11446_/X _11445_/X _11476_/S _15446_/Q sky130_fd_sc_hd__mux2_1
X_14165_ hold545/A _14165_/CLK _14165_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11377_ VGND VPWR VPWR VGND _11377_/X _14846_/Q _11392_/B _14814_/Q sky130_fd_sc_hd__mux2_1
X_10328_ VPWR VGND VPWR VGND _10325_/X _10816_/A _10327_/X _10328_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_1145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10259_ VGND VPWR VGND VPWR _10259_/X _15485_/Q _11003_/A2 _10258_/X _10911_/S sky130_fd_sc_hd__o211a_1
XFILLER_38_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13733__850 VPWR VGND VPWR VGND _15105_/CLK clkload30/A sky130_fd_sc_hd__inv_2
X_14998_ _14998_/Q _14998_/CLK _14998_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_35_833 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_07470_ VPWR VGND VGND VPWR _15448_/Q _07577_/A _07471_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_15619_ _15619_/Q clkload14/A _15619_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09140_ VGND VPWR VPWR VGND _14958_/D clone55/A _09157_/S hold961/X sky130_fd_sc_hd__mux2_1
X_09071_ VGND VPWR VPWR VGND _15022_/D hold1087/X _09090_/S clone55/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08022_ VPWR VGND VGND VPWR _15557_/Q _08022_/B _08023_/B sky130_fd_sc_hd__nor2_1
Xhold701 hold701/X hold701/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold712 hold712/X hold712/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout5 VGND VPWR fanout7/A fanout5/X VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold745 hold745/X hold745/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 hold734/X hold734/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 hold723/X hold723/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ VGND VPWR VGND VPWR _09974_/B _09970_/A _09970_/B _09977_/A _09890_/A sky130_fd_sc_hd__o211a_1
Xhold767 hold767/X hold767/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13582__699 VPWR VGND VPWR VGND _14913_/CLK clkload54/A sky130_fd_sc_hd__inv_2
Xhold778 hold778/X hold778/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 hold756/X hold756/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ VPWR VGND VGND VPWR _08924_/X _15130_/Q _08924_/B sky130_fd_sc_hd__or2_1
Xhold789 hold789/X hold789/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1401 hold1401/X _15321_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1423 hold1423/X _15124_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 hold1412/X _15695_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08855_ VPWR VGND VPWR VGND _08854_/X _15161_/D hold151/X _08853_/Y sky130_fd_sc_hd__a21boi_1
Xhold1434 hold1434/X _14933_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 hold1445/X _15111_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 _07101_/A _15352_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1467 _08914_/A _15135_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_479 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07806_ VGND VPWR VGND VPWR _07809_/A _07868_/A _07867_/A _07867_/B sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08786_ VGND VPWR VPWR VGND _15223_/D _08808_/S fanout76/X hold1146/X sky130_fd_sc_hd__mux2_4
X_07737_ VPWR VGND VPWR VGND _07827_/D _15582_/Q _07714_/X _07739_/B sky130_fd_sc_hd__a21o_1
X_13476__593 VPWR VGND VPWR VGND _14751_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_64_clk _12961__78/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_77_1087 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_685 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07668_ VPWR VGND VGND VPWR _07668_/A _07668_/Y _07668_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_1098 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07599_ VGND VPWR VGND VPWR clone17/A _07421_/A _07561_/X _07599_/X sky130_fd_sc_hd__o21ba_1
X_09407_ VGND VPWR VPWR VGND _14642_/D hold350/X _09414_/S _09826_/A1 sky130_fd_sc_hd__mux2_1
XFILLER_55_1363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09338_ VGND VPWR VPWR VGND _14706_/D hold583/X _09345_/S _09686_/A0 sky130_fd_sc_hd__mux2_1
X_13019__136 VPWR VGND VPWR VGND _14262_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_09269_ VGND VPWR VPWR VGND _14774_/D _09827_/A1 _09269_/S hold605/X sky130_fd_sc_hd__mux2_1
X_11300_ VPWR VGND _14818_/D _11300_/B _11388_/S VPWR VGND sky130_fd_sc_hd__and2_1
X_12919__36 VPWR VGND VPWR VGND _14162_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_12280_ VGND VPWR VPWR VGND _12280_/X hold790/A _12689_/S _14302_/Q sky130_fd_sc_hd__mux2_1
X_11231_ VGND VPWR VPWR VGND _11231_/X _14506_/Q _11231_/S _14186_/Q sky130_fd_sc_hd__mux2_1
X_11162_ VGND VPWR VPWR VGND _11162_/X _11159_/X _11162_/S _11158_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10113_ VGND VPWR VPWR VGND _10113_/X hold626/A _10609_/S hold892/A sky130_fd_sc_hd__mux2_1
X_11093_ VGND VPWR VPWR VGND _11093_/X _14795_/Q _11093_/S _14246_/Q sky130_fd_sc_hd__mux2_1
X_14921_ hold354/A _14921_/CLK _14921_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10044_ VGND VPWR VPWR VGND _10044_/A _15634_/D _10045_/C sky130_fd_sc_hd__xor2_1
XFILLER_75_254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14852_ _14852_/Q clkload26/A _14852_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13717__834 VPWR VGND VPWR VGND _15057_/CLK clkload39/A sky130_fd_sc_hd__inv_2
XFILLER_35_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14783_ hold721/A _14783_/CLK _14783_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11995_ VGND VPWR VPWR VGND _11995_/X _11994_/X _11995_/S _11993_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_55_clk _12936__53/A clkload2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_10946_ VPWR VGND VGND VPWR _10946_/X _11170_/S _10946_/B sky130_fd_sc_hd__or2_1
X_10877_ VGND VPWR VPWR VGND _10877_/X _14368_/Q _11109_/S _14720_/Q sky130_fd_sc_hd__mux2_1
X_15404_ hold315/A _15404_/CLK _15404_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12616_ VPWR VGND VGND VPWR _12616_/X _12624_/S _12616_/B sky130_fd_sc_hd__or2_1
X_15335_ _15335_/Q _15335_/CLK _15335_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12547_ VPWR VGND VGND VPWR _12658_/A _12547_/B _12547_/Y sky130_fd_sc_hd__nor2_1
X_15266_ _15266_/Q _15266_/CLK _15266_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XANTENNA_3 _07593_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_12478_ VGND VPWR VGND VPWR _12478_/X hold729/A _12488_/A2 _12489_/A1 _12477_/X sky130_fd_sc_hd__o211a_1
X_11429_ VGND VPWR VGND VPWR _14929_/D _14930_/Q _11431_/A2 _11428_/X _11431_/C1 sky130_fd_sc_hd__o211a_1
X_15197_ hold201/A _15197_/CLK _15197_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14217_ _14217_/Q _14217_/CLK _14217_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14148_ _14148_/Q _14148_/CLK _14148_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12933__50 VPWR VGND VPWR VGND _14176_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_67_711 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_13163__280 VPWR VGND VPWR VGND _14438_/CLK clkload47/A sky130_fd_sc_hd__inv_2
X_08640_ VPWR VGND VGND VPWR _08640_/X _14392_/Q _08640_/B sky130_fd_sc_hd__or2_1
Xrebuffer26 VPWR VGND VPWR VGND rebuffer26/X rebuffer27/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer15 VPWR VGND VPWR VGND _08233_/A _07564_/B sky130_fd_sc_hd__dlygate4sd1_1
X_14013__1130 VPWR VGND VPWR VGND _15385_/CLK clkload55/A sky130_fd_sc_hd__inv_2
XFILLER_78_1341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08571_ VPWR VGND VGND VPWR _15554_/Q _08571_/Y _08571_/B sky130_fd_sc_hd__nand2_1
Xrebuffer37 VPWR VGND VPWR VGND rebuffer37/X rebuffer38/X sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer48 VPWR VGND VPWR VGND _07883_/B1 _07137_/X sky130_fd_sc_hd__dlygate4sd1_1
Xclkbuf_leaf_46_clk _12970__87/A clkload3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_78_1385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07522_ VGND VPWR VGND VPWR _14803_/Q _14804_/Q _07523_/B sky130_fd_sc_hd__or2_4
X_07453_ VPWR VGND VPWR VGND _15598_/Q _15454_/Q _15599_/Q _07453_/X _15453_/Q sky130_fd_sc_hd__a22o_1
X_07384_ VGND VPWR VPWR VGND _08010_/A _08007_/A _08006_/B _08006_/C sky130_fd_sc_hd__o21ai_4
X_13510__627 VPWR VGND VPWR VGND _14785_/CLK _12961__78/A sky130_fd_sc_hd__inv_2
X_09123_ VGND VPWR VPWR VGND _14972_/D hold433/X _09128_/S _09550_/A1 sky130_fd_sc_hd__mux2_1
X_09054_ VGND VPWR VPWR VGND _15036_/D hold555/X _09059_/S _09688_/A0 sky130_fd_sc_hd__mux2_1
X_08005_ VGND VPWR _08005_/B _08005_/Y _08010_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
Xhold520 hold520/X hold520/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 hold553/X hold553/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 hold542/X hold542/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 hold531/X hold531/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 hold575/X hold575/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 hold586/X hold586/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 hold564/X hold564/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold597/X hold597/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ VGND VPWR VPWR VGND _14126_/D hold1352/X _09956_/S _09955_/X sky130_fd_sc_hd__mux2_1
X_13404__521 VPWR VGND VPWR VGND _14679_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_09887_ VPWR VGND VPWR VGND _09886_/Y _09873_/A _15479_/Q _09887_/X sky130_fd_sc_hd__a21o_1
X_08907_ VGND VPWR VGND VPWR _15139_/D _15138_/Q _08880_/B _08906_/X _11398_/A sky130_fd_sc_hd__o211a_1
Xhold1231 hold1231/X _14795_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 hold1242/X _15340_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ VGND VPWR VPWR VGND _15175_/D fanout17/X _08850_/S hold417/X sky130_fd_sc_hd__mux2_1
Xhold1220 hold1220/X _14790_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 hold1275/X _15434_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 hold1264/X _14837_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 hold1253/X _15157_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 hold1286/X _15334_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 hold1297/X _14842_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ VGND VPWR VPWR VGND _15237_/D fanout9/X _08779_/S hold177/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_clk _12962__79/A clkload5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_54_950 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10800_ VGND VPWR VGND VPWR _10800_/X _10797_/X _10799_/X _11215_/C1 _11218_/A1 sky130_fd_sc_hd__a211o_1
X_11780_ VPWR VGND VGND VPWR _11780_/X hold203/A _12005_/S sky130_fd_sc_hd__or2_1
XFILLER_41_611 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_10731_ VGND VPWR VPWR VGND _10731_/X hold913/A _10743_/B hold418/A sky130_fd_sc_hd__mux2_1
X_14109__1226 VPWR VGND VPWR VGND _15528_/CLK _12923__40/A sky130_fd_sc_hd__inv_2
XFILLER_41_688 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10662_ VGND VPWR VPWR VGND _10662_/X _10661_/X _10662_/S _10660_/X sky130_fd_sc_hd__mux2_1
X_12401_ VGND VPWR VPWR VGND _12401_/X hold843/A _12635_/B hold465/A sky130_fd_sc_hd__mux2_1
X_10593_ VGND VPWR VGND VPWR _10593_/X _10590_/X _10592_/X _10593_/A1 _10741_/C1 sky130_fd_sc_hd__a211o_1
X_15120_ _15120_/Q _15120_/CLK _15120_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12332_ VGND VPWR VGND VPWR _12332_/X _12331_/X _12330_/X _12328_/S _12748_/C1 sky130_fd_sc_hd__a211o_1
X_15051_ hold518/A _15051_/CLK _15051_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12263_ VPWR VGND VGND VPWR _12588_/A1 _12259_/X _12748_/C1 _12263_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_11214_ VPWR VGND VGND VPWR _11214_/X hold329/A _11223_/S sky130_fd_sc_hd__or2_1
XFILLER_64_1429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12194_ VPWR VGND _12194_/X _12193_/X _12189_/X _12176_/S _12185_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_11145_ VGND VPWR VPWR VGND _11145_/X hold930/A _11146_/B hold164/A sky130_fd_sc_hd__mux2_1
X_11076_ VPWR VGND VGND VPWR _11076_/X hold332/A _11186_/S sky130_fd_sc_hd__or2_1
X_13147__264 VPWR VGND VPWR VGND _14422_/CLK clkload12/A sky130_fd_sc_hd__inv_2
XFILLER_7_1345 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14904_ hold356/A _14904_/CLK _14904_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10027_ VPWR VGND _10031_/C _10028_/B _15627_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_49_755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_48_243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_37_917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_23_1148 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14835_ _14835_/Q clkload28/A _14835_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_28_clk clkload45/A clkload4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_5_1080 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14766_ _14766_/Q _14766_/CLK _14766_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11978_ VGND VPWR VPWR VGND _11978_/X hold822/A _12006_/B hold668/A sky130_fd_sc_hd__mux2_1
X_10929_ VGND VPWR VGND VPWR _10929_/X _15021_/Q _12866_/A1 _10928_/X _11244_/S sky130_fd_sc_hd__o211a_1
X_14697_ hold709/A _14697_/CLK _14697_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_75_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13845__962 VPWR VGND VPWR VGND _15217_/CLK _12980__97/A sky130_fd_sc_hd__inv_2
X_15318_ _15318_/Q _15318_/CLK _15318_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13922__1039 VPWR VGND VPWR VGND _15294_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_15249_ _15249_/Q _15249_/CLK _15249_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xfanout329 VGND VPWR _10964_/S _11251_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout318 VPWR VGND _11231_/S _11241_/S VPWR VGND sky130_fd_sc_hd__buf_2
X_09810_ VGND VPWR VPWR VGND _14242_/D fanout57/X _09827_/S hold198/X sky130_fd_sc_hd__mux2_1
Xfanout307 VGND VPWR fanout314/X _10664_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
X_09741_ VGND VPWR VPWR VGND _14305_/D _09757_/S clone46/X hold1170/X sky130_fd_sc_hd__mux2_4
X_09672_ VGND VPWR VPWR VGND _14368_/D _09675_/S hold1222/X fanout50/X sky130_fd_sc_hd__mux2_4
Xclkbuf_leaf_19_clk clkload26/A clkbuf_3_2_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_08623_ VPWR VGND VGND VPWR _08626_/A _08623_/B _08623_/Y sky130_fd_sc_hd__nor2_1
X_08554_ VGND VPWR _08554_/B _08554_/Y _08554_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
X_07505_ VPWR VGND VGND VPWR _15462_/Q _07507_/B _07530_/B sky130_fd_sc_hd__nor2_1
X_08485_ VGND VPWR VGND VPWR _15334_/D hold1193/X _08485_/A2 _08484_/X _08541_/A sky130_fd_sc_hd__o211a_1
XFILLER_51_964 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_1177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07436_ VPWR VGND VGND VPWR _08566_/A _08544_/A _07436_/B sky130_fd_sc_hd__or2_1
X_07367_ VPWR VGND VPWR VGND _07366_/B _07366_/A _10061_/C _08137_/B sky130_fd_sc_hd__a21o_1
XFILLER_6_309 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_09106_ VGND VPWR VPWR VGND _14989_/D hold589/X _09124_/S fanout54/X sky130_fd_sc_hd__mux2_1
X_07298_ VPWR VGND VPWR VGND _07859_/A _07298_/A _07860_/A sky130_fd_sc_hd__or2_2
X_09037_ VGND VPWR VPWR VGND _15053_/D hold688/X _09055_/S fanout54/X sky130_fd_sc_hd__mux2_1
Xhold350 hold350/X hold350/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 hold361/X hold361/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold372/X hold372/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 hold394/X hold394/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/X hold383/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout841 VGND VPWR _12751_/C1 _12677_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout852 VPWR VGND _08277_/S _07966_/A VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout830 VGND VPWR fanout844/X _12085_/C1 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09939_ VGND VPWR VPWR VGND _09937_/Y _09956_/S _09939_/B sky130_fd_sc_hd__and2b_2
Xfanout885 VGND VPWR _07141_/A _10078_/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout863 VPWR VGND _07751_/C _07757_/C VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout874 VGND VPWR _15583_/Q _07119_/A VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xhold1050 hold1050/X _15485_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_405 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_12881_ VPWR VGND VPWR VGND _12878_/C _12883_/A _12878_/A _07421_/A _08195_/A _12878_/B
+ sky130_fd_sc_hd__a2111o_1
Xhold1072 hold1072/X _14868_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 hold1061/X _15488_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 hold1094/X _15003_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ VGND VPWR VPWR VGND _11905_/B hold677/A _12149_/S hold481/A sky130_fd_sc_hd__mux2_1
Xhold1083 hold1083/X _14879_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13788__905 VPWR VGND VPWR VGND _15160_/CLK clkload31/A sky130_fd_sc_hd__inv_2
XFILLER_45_257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11832_ VGND VPWR VGND VPWR _11832_/X _12099_/A1 _11828_/X _11831_/X _12099_/C1 sky130_fd_sc_hd__o211a_1
X_14620_ hold618/A _14620_/CLK _14620_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14551_ hold735/A _14551_/CLK _14551_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11763_ VGND VPWR VPWR VGND _11763_/X _14192_/Q _12086_/S hold404/A sky130_fd_sc_hd__mux2_1
X_13829__946 VPWR VGND VPWR VGND _15201_/CLK clkload53/A sky130_fd_sc_hd__inv_2
X_14482_ hold969/A _14482_/CLK _14482_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11694_ VPWR VGND VPWR VGND _11693_/X _12722_/A1 _11692_/X _11694_/Y sky130_fd_sc_hd__a21oi_1
X_10714_ VGND VPWR VPWR VGND _10714_/X hold682/A _10743_/B hold258/A sky130_fd_sc_hd__mux2_1
X_10645_ VPWR VGND VPWR VGND _10644_/X _10667_/C1 _10643_/X _10645_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_1417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15103_ _15103_/Q _15103_/CLK _15103_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12315_ VPWR VGND VPWR VGND _12314_/X _12596_/C1 _12313_/X _12315_/Y sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_39_Left_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10576_ VPWR VGND VGND VPWR _10576_/X _10732_/S _10576_/B sky130_fd_sc_hd__or2_1
X_12246_ VPWR VGND VGND VPWR _12246_/X hold183/A _12318_/S sky130_fd_sc_hd__or2_1
X_15034_ hold614/A _15034_/CLK _15034_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12903__20 VPWR VGND VPWR VGND _14145_/CLK clkload29/A sky130_fd_sc_hd__inv_2
X_12177_ VPWR VGND VGND VPWR _12214_/A _12177_/B _12177_/Y sky130_fd_sc_hd__nor2_1
X_13381__498 VPWR VGND VPWR VGND _14656_/CLK clkload46/A sky130_fd_sc_hd__inv_2
X_11128_ VGND VPWR VPWR VGND _11128_/X _14279_/Q _11146_/B _14311_/Q sky130_fd_sc_hd__mux2_1
XFILLER_49_541 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_76_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_37_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11059_ VGND VPWR VPWR VGND _11059_/X _11056_/X _11176_/S _11055_/X sky130_fd_sc_hd__mux2_1
X_14818_ _14818_/Q clkload27/A _14818_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_64_599 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14749_ hold508/A _14749_/CLK _14749_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1317 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_783 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08270_ VPWR VGND VGND VPWR _08269_/Y _08172_/X _08270_/A1 _08173_/Y _08270_/X sky130_fd_sc_hd__o22a_1
X_13275__392 VPWR VGND VPWR VGND _14550_/CLK _12955__72/A sky130_fd_sc_hd__inv_2
X_07221_ VPWR VGND _07221_/X _07222_/A _15447_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07152_ VPWR VGND _07154_/A _07153_/B _15475_/Q VPWR VGND sky130_fd_sc_hd__and2_1
X_07083_ VPWR VGND VPWR VGND _09975_/A _10056_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_8_clk clkload14/A clkload0/A VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_13622__739 VPWR VGND VPWR VGND _14962_/CLK clkload47/A sky130_fd_sc_hd__inv_2
Xfanout104 VGND VPWR _08149_/X _09685_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14108__1225 VPWR VGND VPWR VGND _15527_/CLK clkload10/A sky130_fd_sc_hd__inv_2
Xfanout137 VGND VPWR _08730_/B1 _08540_/B1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout126 VGND VPWR _08190_/X _09653_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout115 VGND VPWR _08250_/X _09228_/A0 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xfanout159 VGND VPWR _11421_/X _11439_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout148 VGND VPWR _08686_/A2 _08628_/A2 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_07985_ VGND VPWR VGND VPWR _10074_/A0 _07186_/B _07972_/B _07985_/X _07186_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_09724_ VGND VPWR VPWR VGND _14319_/D _09863_/A0 _09725_/S hold664/X sky130_fd_sc_hd__mux2_1
X_09655_ VGND VPWR VPWR VGND _14415_/D hold839/X _09656_/S _09655_/A0 sky130_fd_sc_hd__mux2_1
X_08606_ VGND VPWR VGND VPWR _08606_/X _08605_/A _08615_/B1 hold1446/X _08605_/Y sky130_fd_sc_hd__a211o_1
Xtt_um_femto_897 uio_out[0] tt_um_femto_897/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xclkbuf_3_2_0_clk clkbuf_3_2_0_clk/X clkbuf_0_clk/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_09586_ VGND VPWR VPWR VGND _14479_/D hold968/X _09587_/S _09863_/A0 sky130_fd_sc_hd__mux2_1
X_13516__633 VPWR VGND VPWR VGND _14791_/CLK clkload41/A sky130_fd_sc_hd__inv_2
X_08537_ VPWR VGND _15318_/D _08537_/B _08541_/A VPWR VGND sky130_fd_sc_hd__and2_1
X_08468_ VPWR VGND VGND VPWR _08468_/X _08468_/A _08482_/B sky130_fd_sc_hd__or2_1
XFILLER_24_975 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07419_ VPWR VGND VGND VPWR _15476_/Q _07145_/X _10074_/A1 _07419_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_1250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08399_ VGND VPWR VPWR VGND _15378_/D fanout17/X _08411_/S hold902/X sky130_fd_sc_hd__mux2_1
X_10430_ VGND VPWR VGND VPWR _10430_/X _10427_/X _10429_/X _10593_/A1 _10667_/C1 sky130_fd_sc_hd__a211o_1
X_10361_ VGND VPWR VPWR VGND _10361_/X hold965/A _10604_/S hold583/A sky130_fd_sc_hd__mux2_1
X_10292_ VGND VPWR VGND VPWR _10292_/X _10291_/X _10290_/X _10510_/S _10630_/C1 sky130_fd_sc_hd__a211o_1
X_12100_ VGND VPWR VPWR VGND _12100_/X _12097_/X _12100_/S _12096_/X sky130_fd_sc_hd__mux2_1
Xhold180 hold180/X hold180/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_12031_ VGND VPWR VPWR VGND _12031_/X _14359_/Q _12043_/B hold502/A sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold191 hold191/X hold191/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout660 _09342_/S _09312_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout682 VGND VPWR _09061_/X _09091_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout693 VPWR VGND _08919_/A2 _08880_/B VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout671 VPWR VGND _09191_/S _09194_/S VPWR VGND sky130_fd_sc_hd__buf_4
X_13921__1038 VPWR VGND VPWR VGND _15293_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_13259__376 VPWR VGND VPWR VGND _14534_/CLK clkload45/A sky130_fd_sc_hd__inv_2
X_12864_ VGND VPWR VPWR VGND _15588_/D _12864_/A1 _14802_/D hold1431/X sky130_fd_sc_hd__mux2_1
XFILLER_27_780 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11815_ VGND VPWR VGND VPWR _11815_/X _12744_/C1 _11810_/X _11814_/X _12864_/A1 sky130_fd_sc_hd__o211a_1
X_12795_ VGND VPWR VGND VPWR _12795_/X _12817_/A _12793_/X _12794_/Y _12807_/A1 sky130_fd_sc_hd__o211a_1
X_15583_ _15583_/Q clkload27/A _15583_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14603_ hold876/A _14603_/CLK _14603_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14534_ _14534_/Q _14534_/CLK _14534_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11746_ VPWR VGND VGND VPWR _11746_/X hold167/A _12409_/B sky130_fd_sc_hd__or2_1
XFILLER_41_271 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_11677_ VPWR VGND VPWR VGND _11676_/X _12029_/A _12195_/B1 _11677_/X sky130_fd_sc_hd__a21o_1
X_14465_ _14465_/Q _14465_/CLK _14465_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10628_ VPWR VGND VGND VPWR _10628_/X hold202/A _10632_/B sky130_fd_sc_hd__or2_1
X_14396_ _14396_/Q clkload18/A _14396_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10559_ VPWR VGND VGND VPWR _10556_/X _10558_/X clone2/A _10559_/X sky130_fd_sc_hd__o21a_1
X_15017_ hold979/A _15017_/CLK _15017_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_12229_ VGND VPWR VGND VPWR _12229_/X _15016_/Q _12229_/A2 _12069_/S _12228_/X sky130_fd_sc_hd__o211a_1
X_07770_ _08256_/B _07766_/Y _07770_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_37_533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13203__320 VPWR VGND VPWR VGND _14478_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_09440_ VGND VPWR VPWR VGND _14612_/D fanout6/X _09441_/S hold677/X sky130_fd_sc_hd__mux2_1
X_09371_ VGND VPWR VPWR VGND _14675_/D hold686/X _09379_/S _09547_/A1 sky130_fd_sc_hd__mux2_1
X_08322_ VGND VPWR VPWR VGND _15497_/D fanout33/X _08330_/S hold909/X sky130_fd_sc_hd__mux2_1
X_12887__4 VPWR VGND VPWR VGND _14129_/CLK clkload25/A sky130_fd_sc_hd__inv_2
X_08253_ VPWR VGND VPWR VGND _08253_/A2 _15334_/Q _08252_/X _08253_/X sky130_fd_sc_hd__a21o_1
X_07204_ VPWR VGND VGND VPWR _08135_/A _08115_/A _07204_/B sky130_fd_sc_hd__or2_1
X_08184_ VPWR VGND VPWR VGND _08180_/A _08280_/A2 _08184_/X _08278_/B _07210_/X _08183_/X
+ sky130_fd_sc_hd__a221o_1
X_07135_ VGND VPWR VGND VPWR _07765_/B _07757_/C _15574_/Q sky130_fd_sc_hd__nand2b_2
X_13052__169 VPWR VGND VPWR VGND _14295_/CLK clkload9/A sky130_fd_sc_hd__inv_2
X_12894__11 VPWR VGND VPWR VGND _14136_/CLK _12891__8/A sky130_fd_sc_hd__inv_2
X_07968_ VPWR VGND VPWR VGND _07345_/C _15461_/Q _07971_/A _07968_/Y sky130_fd_sc_hd__a21oi_1
X_09707_ VGND VPWR VPWR VGND _14336_/D fanout50/X _09725_/S hold973/X sky130_fd_sc_hd__mux2_1
XFILLER_60_1465 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_07899_ VGND VPWR VPWR VGND _07899_/B _07387_/X _07899_/A _07900_/B sky130_fd_sc_hd__or3b_1
XFILLER_21_1449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_823 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09638_ VGND VPWR VPWR VGND _14432_/D hold823/X _09656_/S fanout50/X sky130_fd_sc_hd__mux2_1
XFILLER_3_1381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13750__867 VPWR VGND VPWR VGND _15122_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_09569_ VGND VPWR VPWR VGND _14496_/D hold1016/X _09587_/S _07890_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12580_ VGND VPWR VGND VPWR _12580_/X _12580_/A1 _12576_/X _12579_/X _12702_/C1 sky130_fd_sc_hd__o211a_1
X_11600_ VGND VPWR VGND VPWR _11600_/X hold931/A _12040_/A2 _12008_/A1 _11599_/X sky130_fd_sc_hd__o211a_1
X_11531_ VGND VPWR VPWR VGND _15094_/D _11530_/X _11538_/S _15094_/Q sky130_fd_sc_hd__mux2_1
X_11462_ VGND VPWR VPWR VGND _15071_/D _11461_/X _11480_/S hold1402/X sky130_fd_sc_hd__mux2_1
X_14250_ _14250_/Q _14250_/CLK _14250_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11393_ VGND VPWR VPWR VGND _11393_/X _11418_/S _11393_/S _11368_/A sky130_fd_sc_hd__mux2_1
X_10413_ VPWR VGND _10413_/X _10412_/X _10408_/X clone2/X _10404_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_14181_ hold470/A _14181_/CLK _14181_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10344_ VGND VPWR VPWR VGND _10344_/X hold761/A _10696_/S hold265/A sky130_fd_sc_hd__mux2_1
X_13644__761 VPWR VGND VPWR VGND _14984_/CLK clkload18/A sky130_fd_sc_hd__inv_2
X_10275_ VPWR VGND VPWR VGND _10274_/X _10608_/A1 _10273_/X _10275_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_12014_ VGND VPWR VPWR VGND _12014_/X hold850/A _12112_/S hold187/A sky130_fd_sc_hd__mux2_1
XFILLER_79_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout490 VGND VPWR fanout497/X _11882_/S VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_19_522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_15635_ _15635_/Q clkload49/A _15635_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12847_ VPWR VGND VGND VPWR _12845_/X _12846_/X _11477_/S _15571_/D sky130_fd_sc_hd__o21a_1
X_12778_ VPWR VGND VGND VPWR _12789_/A _08116_/Y _12807_/A1 _12778_/X sky130_fd_sc_hd__o21a_1
X_15566_ _15566_/Q clkload50/A _15566_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_14107__1224 VPWR VGND VPWR VGND _15526_/CLK clkload18/A sky130_fd_sc_hd__inv_2
XFILLER_72_1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14517_ hold180/A _14517_/CLK _14517_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15497_ hold909/A _15497_/CLK _15497_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11729_ VGND VPWR VGND VPWR _11729_/X _12720_/A1 _11725_/X _11728_/X _12485_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_31_1022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_31_1000 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14448_ hold434/A _14448_/CLK _14448_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xhold905 hold905/X hold905/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 hold927/X hold927/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 hold916/X hold916/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ VGND VPWR VGND VPWR _14379_/Q _14379_/D clkload6/A sky130_fd_sc_hd__dfxtp_4
Xhold938 hold938/X hold938/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 hold949/X hold949/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08940_ VPWR VGND VPWR VGND _08969_/A _15126_/Q _08933_/A _08941_/B hold1432/X sky130_fd_sc_hd__a22o_1
X_08871_ VGND VPWR VGND VPWR _15157_/D hold1261/X _08893_/A2 _08870_/X _11315_/A1
+ sky130_fd_sc_hd__o211a_1
X_07822_ VGND VPWR VGND VPWR _07822_/X _07857_/A _07815_/X _07821_/Y _08225_/C1 sky130_fd_sc_hd__o211a_1
X_07753_ VPWR VGND VGND VPWR _07751_/X _07753_/B _08153_/A sky130_fd_sc_hd__nand2b_1
XFILLER_77_1225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07684_ VPWR VGND VPWR VGND _07668_/B _15090_/Q _07881_/A2 _07684_/X _07314_/A sky130_fd_sc_hd__a22o_1
XFILLER_77_1269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09423_ VGND VPWR VPWR VGND _14629_/D fanout69/X _09443_/S hold889/X sky130_fd_sc_hd__mux2_1
XFILLER_53_889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_09354_ VGND VPWR VPWR VGND _14692_/D hold469/X _09357_/S fanout65/X sky130_fd_sc_hd__mux2_1
XFILLER_13_709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08305_ VPWR VGND VPWR VGND _08305_/Y _08318_/S sky130_fd_sc_hd__inv_2
X_13587__704 VPWR VGND VPWR VGND _14918_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
X_09285_ VGND VPWR VPWR VGND _14756_/D fanout66/X _09304_/S hold441/X sky130_fd_sc_hd__mux2_1
X_08236_ VPWR VGND VPWR VGND _08252_/A2 _15156_/Q _08235_/X _08236_/X sky130_fd_sc_hd__a21o_1
X_08167_ VGND VPWR VGND VPWR _08167_/X _08263_/A2 _08164_/X _07206_/X _08166_/X sky130_fd_sc_hd__a211o_1
X_13628__745 VPWR VGND VPWR VGND _14968_/CLK clkload7/A sky130_fd_sc_hd__inv_2
X_07118_ VPWR VGND VPWR VGND _10072_/A _15584_/Q sky130_fd_sc_hd__inv_2
X_13920__1037 VPWR VGND VPWR VGND _15292_/CLK clkload13/A sky130_fd_sc_hd__inv_2
XFILLER_10_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08098_ VPWR VGND VGND VPWR _08147_/A _12781_/A _08098_/Y sky130_fd_sc_hd__nor2_1
X_10060_ VPWR VGND VGND VPWR _10060_/C _14801_/Q _10060_/A _10060_/Y sky130_fd_sc_hd__nor3_1
X_13180__297 VPWR VGND VPWR VGND _14455_/CLK clkload9/A sky130_fd_sc_hd__inv_2
XFILLER_29_897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10962_ VGND VPWR VGND VPWR _10962_/X _15504_/Q _11184_/A2 _10961_/X _11143_/S sky130_fd_sc_hd__o211a_1
X_12701_ VGND VPWR VPWR VGND _12701_/X _14892_/Q _12701_/S hold463/A sky130_fd_sc_hd__mux2_1
XFILLER_70_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10893_ VPWR VGND _10893_/X _10883_/X _10879_/X _12869_/A1 _10893_/B1 VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_44_878 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15420_ hold590/A _15420_/CLK _15420_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12632_ VGND VPWR VGND VPWR _12632_/X _15027_/Q _12743_/A2 _12624_/S _12631_/X sky130_fd_sc_hd__o211a_1
X_15351_ _15351_/Q _15351_/CLK _15351_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12563_ VGND VPWR VGND VPWR _12563_/X _12562_/X _12561_/X _12670_/A1 _12670_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_11_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14302_ _14302_/Q _14302_/CLK _14302_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11514_ VGND VPWR VPWR VGND _11514_/X _15090_/Q _11529_/S _15088_/Q sky130_fd_sc_hd__mux2_1
X_12494_ VGND VPWR VPWR VGND _12494_/X hold900/A _12652_/S hold642/A sky130_fd_sc_hd__mux2_1
X_15282_ hold978/A _15282_/CLK _15282_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13074__191 VPWR VGND VPWR VGND _14317_/CLK clkload24/A sky130_fd_sc_hd__inv_2
X_11445_ VGND VPWR VPWR VGND _11445_/X _15067_/Q _11475_/S _15065_/Q sky130_fd_sc_hd__mux2_1
XFILLER_8_757 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_14233_ hold184/A _14233_/CLK _14233_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11376_ VGND VPWR VPWR VGND _14845_/D _11375_/X _11382_/S hold1307/X sky130_fd_sc_hd__mux2_1
X_14164_ hold453/A _14164_/CLK _14164_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10327_ VPWR VGND VPWR VGND _10326_/X _10851_/A _11259_/C1 _10327_/X sky130_fd_sc_hd__a21o_1
X_10258_ VPWR VGND VGND VPWR _10258_/X hold167/A _10258_/B sky130_fd_sc_hd__or2_1
XFILLER_39_617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_13421__538 VPWR VGND VPWR VGND _14696_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_10189_ VPWR VGND VGND VPWR _10186_/X _10188_/X _10469_/S _10189_/X sky130_fd_sc_hd__o21a_1
X_14997_ hold359/A _14997_/CLK _14997_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_653 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15618_ _15618_/Q clkload27/A _15618_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13315__432 VPWR VGND VPWR VGND _14590_/CLK _12974__91/A sky130_fd_sc_hd__inv_2
X_15549_ _15549_/Q clkload43/A _15549_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_09070_ VGND VPWR VPWR VGND _15023_/D hold1093/X _09091_/S fanout63/X sky130_fd_sc_hd__mux2_1
XFILLER_50_1453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08021_ VPWR VGND VPWR VGND _07426_/X _15620_/Q _08299_/A2 _08032_/A _15584_/Q sky130_fd_sc_hd__a22o_1
XFILLER_11_1437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold702 hold702/X hold702/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 hold735/X hold735/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 hold746/X hold746/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/X hold713/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xfanout6 VPWR VGND fanout6/X fanout7/X VPWR VGND sky130_fd_sc_hd__buf_4
Xhold724 hold724/X hold724/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ VPWR VGND VPWR VGND _08935_/A _07123_/Y _11340_/A _15479_/D sky130_fd_sc_hd__a21oi_1
Xhold757 hold757/X hold757/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 hold779/X hold779/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 hold768/X hold768/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08923_ VGND VPWR VGND VPWR _15131_/D _15130_/Q _08902_/B _08922_/X _08925_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_58_915 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1413 _08939_/B _08938_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08854_ VPWR VGND VGND VPWR hold151/A _08853_/Y _08735_/C _08854_/X sky130_fd_sc_hd__o21a_1
Xhold1402 hold1402/X _15071_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1424 hold1424/X _15080_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1435 hold1435/X _15330_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 hold1446/X _15305_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _08874_/A _15155_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_07805_ VGND VPWR _07888_/B _07710_/A _07868_/A _07888_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_57_458 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1457 hold1457/X _15634_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08785_ VGND VPWR VPWR VGND _15224_/D clone45/X _08808_/S hold171/X sky130_fd_sc_hd__mux2_1
X_07736_ VGND VPWR _07736_/B _08037_/A _07736_/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_37_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07667_ VGND VPWR VGND VPWR _07667_/X _07664_/X _07666_/X _07328_/Y _07333_/Y sky130_fd_sc_hd__a211o_1
XFILLER_0_1373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ VGND VPWR VPWR VGND _14643_/D hold443/X _09406_/S _09859_/A0 sky130_fd_sc_hd__mux2_1
X_07598_ VGND VPWR VPWR VGND _10058_/A1 _07598_/Y _07597_/X _07331_/A sky130_fd_sc_hd__o21ai_4
XFILLER_41_837 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_13058__175 VPWR VGND VPWR VGND _14301_/CLK _12964__81/A sky130_fd_sc_hd__inv_2
X_09337_ VGND VPWR VPWR VGND _14707_/D hold710/X _09345_/S _09685_/A0 sky130_fd_sc_hd__mux2_1
X_09268_ VGND VPWR VPWR VGND _14775_/D _09826_/A1 _09268_/S hold485/X sky130_fd_sc_hd__mux2_1
X_08219_ VPWR VGND VPWR VGND _15545_/Q _15546_/Q _15547_/Q _08220_/C sky130_fd_sc_hd__a21oi_1
X_09199_ VPWR VGND VGND VPWR hold1400/X _09213_/S _09199_/Y sky130_fd_sc_hd__nand2b_1
X_13862__979 VPWR VGND VPWR VGND _15234_/CLK _12951__68/A sky130_fd_sc_hd__inv_2
X_11230_ VGND VPWR VPWR VGND _11234_/B _14634_/Q _11240_/S _14666_/Q sky130_fd_sc_hd__mux2_1
X_11161_ VGND VPWR VGND VPWR _11161_/X _11178_/C1 _11157_/X _11160_/X _11180_/C1 sky130_fd_sc_hd__o211a_1
X_10112_ VGND VPWR VGND VPWR _10112_/X _10109_/X _10111_/X _10614_/A1 _10614_/C1 sky130_fd_sc_hd__a211o_1
XFILLER_76_701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_11092_ VGND VPWR VPWR VGND _11092_/X _11091_/X _11092_/S _11090_/X sky130_fd_sc_hd__mux2_1
X_14106__1223 VPWR VGND VPWR VGND _15525_/CLK clkload13/A sky130_fd_sc_hd__inv_2
X_10043_ VPWR VGND VGND VPWR _10045_/C _10043_/B _15633_/D sky130_fd_sc_hd__nor2_1
X_14920_ hold764/A _14920_/CLK _14920_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13756__873 VPWR VGND VPWR VGND _15128_/CLK _14832_/CLK sky130_fd_sc_hd__inv_2
X_14851_ _14851_/Q clkload26/A _14851_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
X_11994_ VGND VPWR VPWR VGND _11994_/X hold875/A _11998_/S hold870/A sky130_fd_sc_hd__mux2_1
X_14782_ hold384/A _14782_/CLK _14782_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10945_ VGND VPWR VPWR VGND _10945_/X hold716/A _11167_/S hold251/A sky130_fd_sc_hd__mux2_1
X_10876_ VGND VPWR VPWR VGND _10876_/X hold823/A _11109_/S hold697/A sky130_fd_sc_hd__mux2_1
X_12615_ VGND VPWR VPWR VGND _12615_/X hold582/A _12623_/S hold287/A sky130_fd_sc_hd__mux2_1
X_15403_ hold734/A _15403_/CLK _15403_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15334_ _15334_/Q _15334_/CLK _15334_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12546_ VGND VPWR VPWR VGND _12547_/B _12545_/Y _12731_/S _12537_/Y sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_20_Left_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_15265_ _15265_/Q _15265_/CLK _15265_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_12477_ VPWR VGND VGND VPWR _12477_/X hold382/A _12477_/B sky130_fd_sc_hd__or2_1
X_11428_ VGND VPWR VGND VPWR _11428_/X _14929_/Q _11303_/A _11431_/A2 sky130_fd_sc_hd__a21bo_1
XANTENNA_4 _07631_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_15196_ hold186/A _15196_/CLK _15196_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_14216_ _14216_/Q _14216_/CLK _14216_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11359_ VGND VPWR VPWR VGND _11408_/B _11359_/C _11410_/A _11368_/A sky130_fd_sc_hd__or3_2
X_14147_ _14147_/Q _14147_/CLK _14147_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_1413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_08570_ VGND VPWR VGND VPWR _15312_/D hold886/X _08613_/A2 _08569_/X _11337_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_55_929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xrebuffer16 VPWR VGND VPWR VGND _08232_/A _08233_/A sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_54_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xrebuffer27 VPWR VGND VPWR VGND rebuffer27/X rebuffer28/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_48_981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_78_1353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07521_ VPWR VGND VGND VPWR _07534_/B _14803_/Q _14804_/Q sky130_fd_sc_hd__nor2_4
Xrebuffer38 VPWR VGND VPWR VGND rebuffer38/X rebuffer39/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_78_1397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07452_ VPWR VGND VGND VPWR _08575_/A _07452_/B _07496_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_07383_ VGND VPWR VPWR VGND _08025_/A _08006_/C _07381_/X _07379_/X _07258_/B _07088_/Y
+ sky130_fd_sc_hd__a221oi_4
X_09122_ VGND VPWR VPWR VGND _14973_/D hold759/X _09122_/S _09792_/A1 sky130_fd_sc_hd__mux2_1
X_09053_ VGND VPWR VPWR VGND _15037_/D hold495/X _09053_/S _09792_/A1 sky130_fd_sc_hd__mux2_1
X_08004_ VGND VPWR VGND VPWR _07268_/A _08026_/A _08025_/B _08005_/B sky130_fd_sc_hd__o21ba_1
Xhold510 hold510/X hold510/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 hold543/X hold543/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 hold554/X hold554/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_13699__816 VPWR VGND VPWR VGND _15039_/CLK clkload19/A sky130_fd_sc_hd__inv_2
Xhold521 hold521/X hold521/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 hold532/X hold532/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/X hold565/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 hold576/X hold576/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 hold587/X hold587/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ VPWR VGND _09955_/X _09954_/X _09953_/Y _14767_/Q _08492_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_13443__560 VPWR VGND VPWR VGND _14718_/CLK clkload55/A sky130_fd_sc_hd__inv_2
Xhold598 hold598/X hold598/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_09886_ VGND VPWR _09886_/B _09886_/Y _14147_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
X_08906_ VPWR VGND VGND VPWR _08906_/X _15139_/Q _08926_/B sky130_fd_sc_hd__or2_1
XFILLER_58_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1210 hold1210/X _14835_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 hold1221/X _14566_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 hold1232/X _14464_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 _15341_/D _08471_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_08837_ VGND VPWR VPWR VGND _15176_/D _08051_/X _08847_/S hold372/X sky130_fd_sc_hd__mux2_1
Xhold1265 _14837_/D _11350_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 _15158_/D _08869_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 hold1276/X _15148_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_17_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold1287 hold1287/X _15443_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 _14842_/D _11355_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ VGND VPWR VPWR VGND _15238_/D fanout14/X _08779_/S hold232/X sky130_fd_sc_hd__mux2_1
X_07719_ VPWR VGND VPWR VGND _07827_/D _15588_/Q _07714_/X _07721_/B sky130_fd_sc_hd__a21o_1
X_08699_ VGND VPWR VGND VPWR _08699_/X _14392_/Q _08640_/B _08711_/B1 _08639_/X sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_11_Left_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_10730_ VGND VPWR VPWR VGND _10730_/X hold798/A _10730_/S hold722/A sky130_fd_sc_hd__mux2_1
XFILLER_41_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10661_ VGND VPWR VPWR VGND _10661_/X hold918/A _10720_/S hold723/A sky130_fd_sc_hd__mux2_1
X_12400_ VGND VPWR VPWR VGND _12400_/X hold987/A _12409_/B _14689_/Q sky130_fd_sc_hd__mux2_1
X_10592_ VGND VPWR VGND VPWR _10592_/X _15494_/Q _10744_/A2 _10591_/X _10588_/S sky130_fd_sc_hd__o211a_1
X_12331_ VGND VPWR VPWR VGND _12331_/X hold846/A _12339_/B hold786/A sky130_fd_sc_hd__mux2_1
X_12262_ VPWR VGND VGND VPWR _12262_/X _12591_/S _12262_/B sky130_fd_sc_hd__or2_1
X_15050_ hold663/A _15050_/CLK _15050_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11213_ VGND VPWR VPWR VGND _11213_/X _11212_/X _11213_/S _11211_/X sky130_fd_sc_hd__mux2_1
X_12193_ VGND VPWR VGND VPWR _12193_/X _12190_/X _12192_/X _11894_/S _12193_/C1 sky130_fd_sc_hd__a211o_1
X_11144_ VGND VPWR VGND VPWR _11144_/X _11245_/A1 _11143_/X _11140_/X _11255_/C1 sky130_fd_sc_hd__o211a_1
X_11075_ VGND VPWR VPWR VGND _11075_/X hold737/A _11186_/S hold385/A sky130_fd_sc_hd__mux2_1
XFILLER_1_785 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_1324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_10026_ VPWR VGND VGND VPWR _10028_/B _10026_/B _15626_/D sky130_fd_sc_hd__nor2_1
X_14903_ hold644/A _14903_/CLK _14903_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13492__609 VPWR VGND VPWR VGND _14767_/CLK clkload25/A sky130_fd_sc_hd__inv_2
XFILLER_40_1441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_14834_ _14834_/Q clkload29/A _14834_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_29_491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_14765_ _14765_/Q _14765_/CLK _14765_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_11977_ VGND VPWR VPWR VGND _11977_/X hold739/A _12006_/B hold232/A sky130_fd_sc_hd__mux2_1
XFILLER_16_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_10928_ VPWR VGND VGND VPWR _10928_/X hold589/A _11240_/S sky130_fd_sc_hd__or2_1
X_14696_ _14696_/Q _14696_/CLK _14696_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_10859_ VGND VPWR VGND VPWR _14399_/D _12491_/B1 _10857_/X _10858_/X _12677_/C1 sky130_fd_sc_hd__o211a_1
XFILLER_12_380 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15317_ _15317_/Q _15317_/CLK _15317_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13386__503 VPWR VGND VPWR VGND _14661_/CLK _12969__86/A sky130_fd_sc_hd__inv_2
X_12529_ VPWR VGND VGND VPWR _12510_/Y _12528_/X _12677_/A2 _15470_/Q _15470_/D _12677_/C1
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_15248_ hold630/A _15248_/CLK _15248_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_15179_ hold705/A _15179_/CLK _15179_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_13427__544 VPWR VGND VPWR VGND _14702_/CLK _12936__53/A sky130_fd_sc_hd__inv_2
Xfanout308 VGND VPWR _10553_/S _10554_/S VPWR VGND sky130_fd_sc_hd__clkbuf_4
Xfanout319 VGND VPWR _10924_/B _10258_/B VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_09740_ VGND VPWR VPWR VGND _14306_/D fanout58/X _09757_/S hold339/X sky130_fd_sc_hd__mux2_1
.ends

